`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module ZynqAdapter(
  input   clk,
  input   reset,
  output  io_nasti_aw_ready,
  input   io_nasti_aw_valid,
  input  [31:0] io_nasti_aw_bits_addr,
  input  [7:0] io_nasti_aw_bits_len,
  input  [2:0] io_nasti_aw_bits_size,
  input  [1:0] io_nasti_aw_bits_burst,
  input   io_nasti_aw_bits_lock,
  input  [3:0] io_nasti_aw_bits_cache,
  input  [2:0] io_nasti_aw_bits_prot,
  input  [3:0] io_nasti_aw_bits_qos,
  input  [3:0] io_nasti_aw_bits_region,
  input  [11:0] io_nasti_aw_bits_id,
  input   io_nasti_aw_bits_user,
  output  io_nasti_w_ready,
  input   io_nasti_w_valid,
  input  [31:0] io_nasti_w_bits_data,
  input   io_nasti_w_bits_last,
  input  [11:0] io_nasti_w_bits_id,
  input  [3:0] io_nasti_w_bits_strb,
  input   io_nasti_w_bits_user,
  input   io_nasti_b_ready,
  output  io_nasti_b_valid,
  output [1:0] io_nasti_b_bits_resp,
  output [11:0] io_nasti_b_bits_id,
  output  io_nasti_b_bits_user,
  output  io_nasti_ar_ready,
  input   io_nasti_ar_valid,
  input  [31:0] io_nasti_ar_bits_addr,
  input  [7:0] io_nasti_ar_bits_len,
  input  [2:0] io_nasti_ar_bits_size,
  input  [1:0] io_nasti_ar_bits_burst,
  input   io_nasti_ar_bits_lock,
  input  [3:0] io_nasti_ar_bits_cache,
  input  [2:0] io_nasti_ar_bits_prot,
  input  [3:0] io_nasti_ar_bits_qos,
  input  [3:0] io_nasti_ar_bits_region,
  input  [11:0] io_nasti_ar_bits_id,
  input   io_nasti_ar_bits_user,
  input   io_nasti_r_ready,
  output  io_nasti_r_valid,
  output [1:0] io_nasti_r_bits_resp,
  output [31:0] io_nasti_r_bits_data,
  output  io_nasti_r_bits_last,
  output [11:0] io_nasti_r_bits_id,
  output  io_nasti_r_bits_user,
  output  io_reset,
  input   io_debug_req_ready,
  output  io_debug_req_valid,
  output [4:0] io_debug_req_bits_addr,
  output [33:0] io_debug_req_bits_data,
  output [1:0] io_debug_req_bits_op,
  output  io_debug_resp_ready,
  input   io_debug_resp_valid,
  input  [33:0] io_debug_resp_bits_data,
  input  [1:0] io_debug_resp_bits_resp
);
  wire  T_371_valid;
  wire [4:0] T_371_bits_addr;
  wire [33:0] T_371_bits_data;
  wire [1:0] T_371_bits_op;
  reg  reqReg_valid;
  reg [31:0] GEN_39;
  reg [4:0] reqReg_bits_addr;
  reg [31:0] GEN_40;
  reg [33:0] reqReg_bits_data;
  reg [63:0] GEN_41;
  reg [1:0] reqReg_bits_op;
  reg [31:0] GEN_42;
  wire  T_402_valid;
  wire [33:0] T_402_bits_data;
  wire [1:0] T_402_bits_resp;
  reg  respReg_valid;
  reg [31:0] GEN_43;
  reg [33:0] respReg_bits_data;
  reg [63:0] GEN_44;
  reg [1:0] respReg_bits_resp;
  reg [31:0] GEN_45;
  wire  T_420;
  reg  awReady;
  reg [31:0] GEN_46;
  wire  GEN_0;
  wire  T_423;
  wire  T_424;
  reg  wReady;
  reg [31:0] GEN_47;
  wire  GEN_1;
  reg  arReady;
  reg [31:0] GEN_48;
  reg  rValid;
  reg [31:0] GEN_49;
  reg  bValid;
  reg [31:0] GEN_50;
  reg [11:0] bId;
  reg [31:0] GEN_51;
  wire [11:0] GEN_2;
  wire  T_429;
  reg [11:0] rId;
  reg [31:0] GEN_52;
  wire [11:0] GEN_3;
  reg [31:0] wData;
  reg [31:0] GEN_53;
  wire [31:0] GEN_4;
  wire [5:0] T_432;
  reg [5:0] wAddr;
  reg [31:0] GEN_54;
  wire [5:0] GEN_5;
  wire [5:0] T_434;
  reg [5:0] rAddr;
  reg [31:0] GEN_55;
  wire [5:0] GEN_6;
  reg  resetReg;
  reg [31:0] GEN_56;
  wire  T_437;
  wire [1:0] T_438;
  wire [3:0] T_439;
  wire [31:0] T_440;
  wire [31:0] rData;
  wire  T_443;
  wire  T_444;
  wire  T_447;
  wire  T_448;
  wire  T_449;
  wire  GEN_7;
  wire  T_451;
  wire  T_453;
  wire  GEN_8;
  wire  GEN_9;
  wire  T_457;
  wire  T_459;
  wire  T_460;
  wire  GEN_10;
  wire  T_465;
  wire  T_466;
  wire  T_467;
  wire [4:0] T_468;
  wire [1:0] T_469;
  wire [1:0] T_470;
  wire [31:0] T_471;
  wire [33:0] T_472;
  wire [4:0] GEN_11;
  wire [1:0] GEN_12;
  wire [33:0] GEN_13;
  wire  T_474;
  wire [1:0] T_475;
  wire [33:0] T_476;
  wire [33:0] GEN_14;
  wire [4:0] GEN_15;
  wire [1:0] GEN_16;
  wire [33:0] GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [4:0] GEN_21;
  wire [1:0] GEN_22;
  wire [33:0] GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  T_482;
  wire  T_483;
  wire  GEN_28;
  wire  T_485;
  wire  GEN_29;
  wire  T_487;
  wire  GEN_30;
  wire [33:0] GEN_31;
  wire [1:0] GEN_32;
  wire  GEN_33;
  wire [1:0] T_498_resp;
  wire [31:0] T_498_data;
  wire  T_498_last;
  wire [11:0] T_498_id;
  wire  T_498_user;
  wire [1:0] T_510_resp;
  wire [11:0] T_510_id;
  wire  T_510_user;
  wire  T_515;
  wire  T_517;
  wire [3:0] T_518;
  wire  T_520;
  wire  T_521;
  wire  T_522;
  wire  T_524;
  wire  T_526;
  wire  T_528;
  wire  T_529;
  wire  T_537;
  wire  T_538;
  wire  T_539;
  wire  T_541;
  wire  T_543;
  wire  T_545;
  wire  T_546;
  wire  T_547;
  wire  T_548;
  wire  T_549;
  wire  T_551;
  wire [4:0] GEN_34;
  reg [31:0] GEN_57;
  wire [33:0] GEN_35;
  reg [63:0] GEN_58;
  wire [1:0] GEN_36;
  reg [31:0] GEN_59;
  wire [33:0] GEN_37;
  reg [63:0] GEN_60;
  wire [1:0] GEN_38;
  reg [31:0] GEN_61;
  assign io_nasti_aw_ready = awReady;
  assign io_nasti_w_ready = wReady;
  assign io_nasti_b_valid = bValid;
  assign io_nasti_b_bits_resp = T_510_resp;
  assign io_nasti_b_bits_id = T_510_id;
  assign io_nasti_b_bits_user = T_510_user;
  assign io_nasti_ar_ready = respReg_valid;
  assign io_nasti_r_valid = rValid;
  assign io_nasti_r_bits_resp = T_498_resp;
  assign io_nasti_r_bits_data = T_498_data;
  assign io_nasti_r_bits_last = T_498_last;
  assign io_nasti_r_bits_id = T_498_id;
  assign io_nasti_r_bits_user = T_498_user;
  assign io_reset = resetReg;
  assign io_debug_req_valid = reqReg_valid;
  assign io_debug_req_bits_addr = reqReg_bits_addr;
  assign io_debug_req_bits_data = reqReg_bits_data;
  assign io_debug_req_bits_op = reqReg_bits_op;
  assign io_debug_resp_ready = T_515;
  assign T_371_valid = 1'h0;
  assign T_371_bits_addr = GEN_34;
  assign T_371_bits_data = GEN_35;
  assign T_371_bits_op = GEN_36;
  assign T_402_valid = 1'h0;
  assign T_402_bits_data = GEN_37;
  assign T_402_bits_resp = GEN_38;
  assign T_420 = io_nasti_aw_ready & io_nasti_aw_valid;
  assign GEN_0 = T_420 ? 1'h0 : awReady;
  assign T_423 = io_nasti_w_ready & io_nasti_w_valid;
  assign T_424 = T_423 & io_nasti_w_bits_last;
  assign GEN_1 = T_424 ? 1'h0 : wReady;
  assign GEN_2 = T_420 ? io_nasti_aw_bits_id : bId;
  assign T_429 = io_nasti_ar_ready & io_nasti_ar_valid;
  assign GEN_3 = T_429 ? io_nasti_ar_bits_id : rId;
  assign GEN_4 = T_424 ? io_nasti_w_bits_data : wData;
  assign T_432 = io_nasti_aw_bits_addr[5:0];
  assign GEN_5 = T_420 ? T_432 : wAddr;
  assign T_434 = io_nasti_ar_bits_addr[5:0];
  assign GEN_6 = T_429 ? T_434 : rAddr;
  assign T_437 = rAddr[2];
  assign T_438 = respReg_bits_data[33:32];
  assign T_439 = {respReg_bits_resp,T_438};
  assign T_440 = respReg_bits_data[31:0];
  assign rData = T_437 ? {{28'd0}, T_439} : T_440;
  assign T_443 = ~ io_nasti_aw_ready;
  assign T_444 = T_420 | T_443;
  assign T_447 = ~ io_nasti_w_ready;
  assign T_448 = T_424 | T_447;
  assign T_449 = T_444 & T_448;
  assign GEN_7 = T_449 ? 1'h1 : bValid;
  assign T_451 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_453 = wAddr == 6'h8;
  assign GEN_8 = T_453 ? 1'h1 : reqReg_valid;
  assign GEN_9 = T_453 ? 1'h0 : respReg_valid;
  assign T_457 = wAddr == 6'h20;
  assign T_459 = T_453 == 1'h0;
  assign T_460 = T_459 & T_457;
  assign GEN_10 = T_460 ? 1'h1 : resetReg;
  assign T_465 = T_457 == 1'h0;
  assign T_466 = T_459 & T_465;
  assign T_467 = wAddr[2];
  assign T_468 = wData[8:4];
  assign T_469 = wData[3:2];
  assign T_470 = wData[1:0];
  assign T_471 = reqReg_bits_data[31:0];
  assign T_472 = {T_470,T_471};
  assign GEN_11 = T_467 ? T_468 : reqReg_bits_addr;
  assign GEN_12 = T_467 ? T_469 : reqReg_bits_op;
  assign GEN_13 = T_467 ? T_472 : reqReg_bits_data;
  assign T_474 = T_467 == 1'h0;
  assign T_475 = reqReg_bits_data[33:32];
  assign T_476 = {T_475,wData};
  assign GEN_14 = T_474 ? T_476 : GEN_13;
  assign GEN_15 = T_466 ? GEN_11 : reqReg_bits_addr;
  assign GEN_16 = T_466 ? GEN_12 : reqReg_bits_op;
  assign GEN_17 = T_466 ? GEN_14 : reqReg_bits_data;
  assign GEN_18 = T_451 ? GEN_8 : reqReg_valid;
  assign GEN_19 = T_451 ? GEN_9 : respReg_valid;
  assign GEN_20 = T_451 ? GEN_10 : resetReg;
  assign GEN_21 = T_451 ? GEN_15 : reqReg_bits_addr;
  assign GEN_22 = T_451 ? GEN_16 : reqReg_bits_op;
  assign GEN_23 = T_451 ? GEN_17 : reqReg_bits_data;
  assign GEN_24 = T_451 ? 1'h1 : GEN_0;
  assign GEN_25 = T_451 ? 1'h1 : GEN_1;
  assign GEN_26 = T_451 ? 1'h0 : GEN_7;
  assign GEN_27 = T_429 ? 1'h1 : rValid;
  assign T_482 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_483 = T_482 & io_nasti_r_bits_last;
  assign GEN_28 = T_483 ? 1'h0 : GEN_27;
  assign T_485 = io_debug_req_ready & io_debug_req_valid;
  assign GEN_29 = T_485 ? 1'h0 : GEN_18;
  assign T_487 = io_debug_resp_ready & io_debug_resp_valid;
  assign GEN_30 = T_487 ? 1'h1 : GEN_19;
  assign GEN_31 = T_487 ? io_debug_resp_bits_data : respReg_bits_data;
  assign GEN_32 = T_487 ? io_debug_resp_bits_resp : respReg_bits_resp;
  assign GEN_33 = resetReg ? 1'h0 : GEN_20;
  assign T_498_resp = 2'h0;
  assign T_498_data = rData;
  assign T_498_last = 1'h1;
  assign T_498_id = rId;
  assign T_498_user = 1'h0;
  assign T_510_resp = 2'h0;
  assign T_510_id = bId;
  assign T_510_user = 1'h0;
  assign T_515 = ~ respReg_valid;
  assign T_517 = io_nasti_w_valid == 1'h0;
  assign T_518 = ~ io_nasti_w_bits_strb;
  assign T_520 = T_518 == 4'h0;
  assign T_521 = T_517 | T_520;
  assign T_522 = T_521 | reset;
  assign T_524 = T_522 == 1'h0;
  assign T_526 = io_nasti_ar_valid == 1'h0;
  assign T_528 = io_nasti_ar_bits_len == 8'h0;
  assign T_529 = T_526 | T_528;
  assign T_537 = io_nasti_ar_bits_burst == 2'h0;
  assign T_538 = T_529 | T_537;
  assign T_539 = T_538 | reset;
  assign T_541 = T_539 == 1'h0;
  assign T_543 = io_nasti_aw_valid == 1'h0;
  assign T_545 = io_nasti_aw_bits_len == 8'h0;
  assign T_546 = T_543 | T_545;
  assign T_547 = io_nasti_aw_bits_burst == 2'h0;
  assign T_548 = T_546 | T_547;
  assign T_549 = T_548 | reset;
  assign T_551 = T_549 == 1'h0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_34 = GEN_57[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_35 = GEN_58[33:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_36 = GEN_59[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_37 = GEN_60[33:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_38 = GEN_61[1:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  reqReg_valid = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  reqReg_bits_addr = GEN_40[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {2{$random}};
  reqReg_bits_data = GEN_41[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  reqReg_bits_op = GEN_42[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  respReg_valid = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {2{$random}};
  respReg_bits_data = GEN_44[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  respReg_bits_resp = GEN_45[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_46 = {1{$random}};
  awReady = GEN_46[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  wReady = GEN_47[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  arReady = GEN_48[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_49 = {1{$random}};
  rValid = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  bValid = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {1{$random}};
  bId = GEN_51[11:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  rId = GEN_52[11:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {1{$random}};
  wData = GEN_53[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {1{$random}};
  wAddr = GEN_54[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {1{$random}};
  rAddr = GEN_55[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {1{$random}};
  resetReg = GEN_56[0:0];
  `endif
  GEN_57 = {1{$random}};
  GEN_58 = {2{$random}};
  GEN_59 = {1{$random}};
  GEN_60 = {2{$random}};
  GEN_61 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      reqReg_valid <= T_371_valid;
    end else begin
      if(T_485) begin
        reqReg_valid <= 1'h0;
      end else begin
        if(T_451) begin
          if(T_453) begin
            reqReg_valid <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      reqReg_bits_addr <= T_371_bits_addr;
    end else begin
      if(T_451) begin
        if(T_466) begin
          if(T_467) begin
            reqReg_bits_addr <= T_468;
          end
        end
      end
    end
    if(reset) begin
      reqReg_bits_data <= T_371_bits_data;
    end else begin
      if(T_451) begin
        if(T_466) begin
          if(T_474) begin
            reqReg_bits_data <= T_476;
          end else begin
            if(T_467) begin
              reqReg_bits_data <= T_472;
            end
          end
        end
      end
    end
    if(reset) begin
      reqReg_bits_op <= T_371_bits_op;
    end else begin
      if(T_451) begin
        if(T_466) begin
          if(T_467) begin
            reqReg_bits_op <= T_469;
          end
        end
      end
    end
    if(reset) begin
      respReg_valid <= T_402_valid;
    end else begin
      if(T_487) begin
        respReg_valid <= 1'h1;
      end else begin
        if(T_451) begin
          if(T_453) begin
            respReg_valid <= 1'h0;
          end
        end
      end
    end
    if(reset) begin
      respReg_bits_data <= T_402_bits_data;
    end else begin
      if(T_487) begin
        respReg_bits_data <= io_debug_resp_bits_data;
      end
    end
    if(reset) begin
      respReg_bits_resp <= T_402_bits_resp;
    end else begin
      if(T_487) begin
        respReg_bits_resp <= io_debug_resp_bits_resp;
      end
    end
    if(reset) begin
      awReady <= 1'h1;
    end else begin
      if(T_451) begin
        awReady <= 1'h1;
      end else begin
        if(T_420) begin
          awReady <= 1'h0;
        end
      end
    end
    if(reset) begin
      wReady <= 1'h1;
    end else begin
      if(T_451) begin
        wReady <= 1'h1;
      end else begin
        if(T_424) begin
          wReady <= 1'h0;
        end
      end
    end
    if(reset) begin
      arReady <= 1'h0;
    end
    if(reset) begin
      rValid <= 1'h0;
    end else begin
      if(T_483) begin
        rValid <= 1'h0;
      end else begin
        if(T_429) begin
          rValid <= 1'h1;
        end
      end
    end
    if(reset) begin
      bValid <= 1'h0;
    end else begin
      if(T_451) begin
        bValid <= 1'h0;
      end else begin
        if(T_449) begin
          bValid <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_420) begin
        bId <= io_nasti_aw_bits_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_429) begin
        rId <= io_nasti_ar_bits_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_424) begin
        wData <= io_nasti_w_bits_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_420) begin
        wAddr <= T_432;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_429) begin
        rAddr <= T_434;
      end
    end
    if(reset) begin
      resetReg <= 1'h0;
    end else begin
      if(resetReg) begin
        resetReg <= 1'h0;
      end else begin
        if(T_451) begin
          if(T_460) begin
            resetReg <= 1'h1;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_524) begin
          $fwrite(32'h80000002,"Assertion failed: Nasti to DebugBusIO converter cannot take partial writes\n    at Adapter.scala:129 assert(!w.valid || w.bits.strb.andR,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_524) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_541) begin
          $fwrite(32'h80000002,"Assertion failed: Nasti to DebugBusIO converter can only take fixed bursts\n    at Adapter.scala:131 assert(!ar.valid ||\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_541) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_551) begin
          $fwrite(32'h80000002,"Assertion failed: Nasti to DebugBusIO converter can only take fixed bursts\n    at Adapter.scala:135 assert(!aw.valid ||\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_551) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module RVCExpander(
  input   clk,
  input   reset,
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0] io_out_rd,
  output [4:0] io_out_rs1,
  output [4:0] io_out_rs2,
  output [4:0] io_out_rs3,
  output  io_rvc
);
  wire [1:0] T_8;
  wire  T_10;
  wire [7:0] T_11;
  wire  T_13;
  wire [6:0] T_16;
  wire [3:0] T_17;
  wire [1:0] T_18;
  wire  T_19;
  wire  T_20;
  wire [2:0] T_22;
  wire [5:0] T_23;
  wire [6:0] T_24;
  wire [9:0] T_25;
  wire [2:0] T_29;
  wire [4:0] T_30;
  wire [11:0] T_31;
  wire [14:0] T_32;
  wire [17:0] T_33;
  wire [29:0] T_34;
  wire [4:0] T_42;
  wire [31:0] T_49_bits;
  wire [4:0] T_49_rd;
  wire [4:0] T_49_rs1;
  wire [4:0] T_49_rs2;
  wire [4:0] T_49_rs3;
  wire [1:0] T_55;
  wire [2:0] T_56;
  wire [4:0] T_58;
  wire [7:0] T_59;
  wire [2:0] T_61;
  wire [4:0] T_62;
  wire [11:0] T_68;
  wire [12:0] T_69;
  wire [15:0] T_70;
  wire [27:0] T_71;
  wire [31:0] T_88_bits;
  wire [4:0] T_88_rd;
  wire [4:0] T_88_rs1;
  wire [4:0] T_88_rs2;
  wire [4:0] T_88_rs3;
  wire [3:0] T_99;
  wire [6:0] T_100;
  wire [11:0] T_109;
  wire [11:0] T_110;
  wire [14:0] T_111;
  wire [26:0] T_112;
  wire [31:0] T_129_bits;
  wire [4:0] T_129_rd;
  wire [4:0] T_129_rs1;
  wire [4:0] T_129_rs2;
  wire [4:0] T_129_rs3;
  wire [27:0] T_151;
  wire [31:0] T_168_bits;
  wire [4:0] T_168_rd;
  wire [4:0] T_168_rs1;
  wire [4:0] T_168_rs2;
  wire [4:0] T_168_rs3;
  wire [1:0] T_181;
  wire [4:0] T_196;
  wire [7:0] T_198;
  wire [14:0] T_199;
  wire [6:0] T_200;
  wire [11:0] T_201;
  wire [26:0] T_202;
  wire [31:0] T_219_bits;
  wire [4:0] T_219_rd;
  wire [4:0] T_219_rs1;
  wire [4:0] T_219_rs2;
  wire [4:0] T_219_rs3;
  wire [2:0] T_230;
  wire [4:0] T_243;
  wire [7:0] T_245;
  wire [14:0] T_246;
  wire [7:0] T_247;
  wire [12:0] T_248;
  wire [27:0] T_249;
  wire [31:0] T_266_bits;
  wire [4:0] T_266_rd;
  wire [4:0] T_266_rs1;
  wire [4:0] T_266_rs2;
  wire [4:0] T_266_rs3;
  wire [14:0] T_297;
  wire [26:0] T_300;
  wire [31:0] T_317_bits;
  wire [4:0] T_317_rd;
  wire [4:0] T_317_rs1;
  wire [4:0] T_317_rs2;
  wire [4:0] T_317_rs3;
  wire [14:0] T_344;
  wire [27:0] T_347;
  wire [31:0] T_364_bits;
  wire [4:0] T_364_rd;
  wire [4:0] T_364_rs1;
  wire [4:0] T_364_rs2;
  wire [4:0] T_364_rs3;
  wire  T_370;
  wire [6:0] T_374;
  wire [4:0] T_375;
  wire [11:0] T_376;
  wire [4:0] T_377;
  wire [11:0] T_381;
  wire [16:0] T_382;
  wire [19:0] T_383;
  wire [31:0] T_384;
  wire [31:0] T_397_bits;
  wire [4:0] T_397_rd;
  wire [4:0] T_397_rs1;
  wire [4:0] T_397_rs2;
  wire [4:0] T_397_rs3;
  wire  T_405;
  wire [6:0] T_408;
  wire [11:0] T_419;
  wire [31:0] T_422;
  wire [31:0] T_435_bits;
  wire [4:0] T_435_rd;
  wire [4:0] T_435_rs1;
  wire [4:0] T_435_rs2;
  wire [4:0] T_435_rs3;
  wire [16:0] T_453;
  wire [19:0] T_454;
  wire [31:0] T_455;
  wire [31:0] T_468_bits;
  wire [4:0] T_468_rd;
  wire [4:0] T_468_rs1;
  wire [4:0] T_468_rs2;
  wire [4:0] T_468_rs3;
  wire  T_482;
  wire [6:0] T_485;
  wire [14:0] T_490;
  wire [19:0] T_493;
  wire [31:0] T_494;
  wire [19:0] T_495;
  wire [24:0] T_497;
  wire [31:0] T_498;
  wire [31:0] T_511_bits;
  wire [4:0] T_511_rd;
  wire [4:0] T_511_rs1;
  wire [4:0] T_511_rs2;
  wire [4:0] T_511_rs3;
  wire  T_519;
  wire  T_522;
  wire  T_523;
  wire [6:0] T_535;
  wire [2:0] T_540;
  wire [1:0] T_541;
  wire  T_543;
  wire [1:0] T_546;
  wire [5:0] T_547;
  wire [4:0] T_548;
  wire [5:0] T_549;
  wire [11:0] T_550;
  wire [11:0] T_554;
  wire [16:0] T_555;
  wire [19:0] T_556;
  wire [31:0] T_557;
  wire [31:0] T_570_bits;
  wire [4:0] T_570_rd;
  wire [4:0] T_570_rs1;
  wire [4:0] T_570_rs2;
  wire [4:0] T_570_rs3;
  wire [31:0] T_576_bits;
  wire [4:0] T_576_rd;
  wire [4:0] T_576_rs1;
  wire [4:0] T_576_rs2;
  wire [4:0] T_576_rs3;
  wire [5:0] T_584;
  wire [11:0] T_593;
  wire [10:0] T_594;
  wire [13:0] T_595;
  wire [25:0] T_596;
  wire [30:0] GEN_0;
  wire [30:0] T_613;
  wire [16:0] T_630;
  wire [19:0] T_631;
  wire [31:0] T_632;
  wire [2:0] T_643;
  wire [2:0] T_645;
  wire  T_647;
  wire [2:0] T_649;
  wire  T_651;
  wire  T_655;
  wire [1:0] T_656;
  wire [1:0] T_662;
  wire [2:0] T_671;
  wire [2:0] T_676;
  wire [2:0] T_677;
  wire [2:0] T_678;
  wire  T_681;
  wire [30:0] T_684;
  wire [6:0] T_688;
  wire [11:0] T_698;
  wire [9:0] T_699;
  wire [12:0] T_700;
  wire [24:0] T_701;
  wire [30:0] GEN_1;
  wire [30:0] T_702;
  wire [1:0] T_703;
  wire [1:0] T_705;
  wire  T_707;
  wire  T_711;
  wire [31:0] T_712;
  wire [30:0] T_717;
  wire [31:0] T_718;
  wire [31:0] T_735_bits;
  wire [4:0] T_735_rd;
  wire [4:0] T_735_rs1;
  wire [4:0] T_735_rs2;
  wire [4:0] T_735_rs3;
  wire [9:0] T_745;
  wire  T_746;
  wire [1:0] T_747;
  wire  T_749;
  wire  T_751;
  wire [2:0] T_752;
  wire [3:0] T_754;
  wire [1:0] T_755;
  wire [5:0] T_756;
  wire [1:0] T_757;
  wire [10:0] T_758;
  wire [12:0] T_759;
  wire [14:0] T_760;
  wire [20:0] T_761;
  wire  T_762;
  wire [9:0] T_784;
  wire  T_806;
  wire [7:0] T_828;
  wire [12:0] T_831;
  wire [19:0] T_832;
  wire [10:0] T_833;
  wire [11:0] T_834;
  wire [31:0] T_835;
  wire [31:0] T_850_bits;
  wire [4:0] T_850_rd;
  wire [4:0] T_850_rs1;
  wire [4:0] T_850_rs2;
  wire [4:0] T_850_rs3;
  wire [4:0] T_860;
  wire [3:0] T_866;
  wire [4:0] T_867;
  wire [6:0] T_868;
  wire [7:0] T_869;
  wire [12:0] T_870;
  wire  T_871;
  wire [5:0] T_887;
  wire [3:0] T_908;
  wire  T_924;
  wire [7:0] T_926;
  wire [6:0] T_927;
  wire [14:0] T_928;
  wire [9:0] T_929;
  wire [6:0] T_930;
  wire [16:0] T_931;
  wire [31:0] T_932;
  wire [31:0] T_947_bits;
  wire [4:0] T_947_rd;
  wire [4:0] T_947_rs1;
  wire [4:0] T_947_rs2;
  wire [4:0] T_947_rs3;
  wire [6:0] T_1024;
  wire [14:0] T_1025;
  wire [31:0] T_1029;
  wire [31:0] T_1042_bits;
  wire [4:0] T_1042_rd;
  wire [4:0] T_1042_rs1;
  wire [4:0] T_1042_rs2;
  wire [4:0] T_1042_rs3;
  wire [10:0] T_1056;
  wire [13:0] T_1057;
  wire [25:0] T_1058;
  wire [31:0] T_1069_bits;
  wire [4:0] T_1069_rd;
  wire [4:0] T_1069_rs1;
  wire [4:0] T_1069_rs2;
  wire [4:0] T_1069_rs3;
  wire [4:0] T_1079;
  wire [3:0] T_1080;
  wire [8:0] T_1081;
  wire [11:0] T_1086;
  wire [13:0] T_1087;
  wire [16:0] T_1088;
  wire [28:0] T_1089;
  wire [31:0] T_1100_bits;
  wire [4:0] T_1100_rd;
  wire [4:0] T_1100_rs1;
  wire [4:0] T_1100_rs2;
  wire [4:0] T_1100_rs3;
  wire [1:0] T_1106;
  wire [2:0] T_1108;
  wire [4:0] T_1110;
  wire [2:0] T_1111;
  wire [7:0] T_1112;
  wire [11:0] T_1117;
  wire [12:0] T_1118;
  wire [15:0] T_1119;
  wire [27:0] T_1120;
  wire [31:0] T_1131_bits;
  wire [4:0] T_1131_rd;
  wire [4:0] T_1131_rs1;
  wire [4:0] T_1131_rs2;
  wire [4:0] T_1131_rs3;
  wire [28:0] T_1151;
  wire [31:0] T_1162_bits;
  wire [4:0] T_1162_rd;
  wire [4:0] T_1162_rs1;
  wire [4:0] T_1162_rs2;
  wire [4:0] T_1162_rs3;
  wire [11:0] T_1173;
  wire [9:0] T_1174;
  wire [12:0] T_1175;
  wire [24:0] T_1176;
  wire [31:0] T_1187_bits;
  wire [4:0] T_1187_rd;
  wire [4:0] T_1187_rs1;
  wire [4:0] T_1187_rs2;
  wire [4:0] T_1187_rs3;
  wire [9:0] T_1199;
  wire [12:0] T_1200;
  wire [24:0] T_1201;
  wire [31:0] T_1212_bits;
  wire [4:0] T_1212_rd;
  wire [4:0] T_1212_rs1;
  wire [4:0] T_1212_rs2;
  wire [4:0] T_1212_rs3;
  wire [24:0] T_1226;
  wire [17:0] T_1227;
  wire [24:0] T_1229;
  wire [24:0] T_1233;
  wire [31:0] T_1244_bits;
  wire [4:0] T_1244_rd;
  wire [4:0] T_1244_rs1;
  wire [4:0] T_1244_rs2;
  wire [4:0] T_1244_rs3;
  wire  T_1252;
  wire [31:0] T_1253_bits;
  wire [4:0] T_1253_rd;
  wire [4:0] T_1253_rs1;
  wire [4:0] T_1253_rs2;
  wire [4:0] T_1253_rs3;
  wire [24:0] T_1267;
  wire [24:0] T_1270;
  wire [24:0] T_1272;
  wire [24:0] T_1276;
  wire [31:0] T_1287_bits;
  wire [4:0] T_1287_rd;
  wire [4:0] T_1287_rs1;
  wire [4:0] T_1287_rs2;
  wire [4:0] T_1287_rs3;
  wire [31:0] T_1296_bits;
  wire [4:0] T_1296_rd;
  wire [4:0] T_1296_rs1;
  wire [4:0] T_1296_rs2;
  wire [4:0] T_1296_rs3;
  wire [31:0] T_1303_bits;
  wire [4:0] T_1303_rd;
  wire [4:0] T_1303_rs1;
  wire [4:0] T_1303_rs2;
  wire [4:0] T_1303_rs3;
  wire [5:0] T_1312;
  wire [8:0] T_1313;
  wire [3:0] T_1314;
  wire [4:0] T_1323;
  wire [7:0] T_1325;
  wire [14:0] T_1326;
  wire [8:0] T_1327;
  wire [13:0] T_1328;
  wire [28:0] T_1329;
  wire [31:0] T_1340_bits;
  wire [4:0] T_1340_rd;
  wire [4:0] T_1340_rs1;
  wire [4:0] T_1340_rs2;
  wire [4:0] T_1340_rs3;
  wire [1:0] T_1346;
  wire [3:0] T_1347;
  wire [5:0] T_1349;
  wire [7:0] T_1350;
  wire [2:0] T_1351;
  wire [4:0] T_1360;
  wire [7:0] T_1362;
  wire [14:0] T_1363;
  wire [7:0] T_1364;
  wire [12:0] T_1365;
  wire [27:0] T_1366;
  wire [31:0] T_1377_bits;
  wire [4:0] T_1377_rd;
  wire [4:0] T_1377_rs1;
  wire [4:0] T_1377_rs2;
  wire [4:0] T_1377_rs3;
  wire [14:0] T_1400;
  wire [28:0] T_1403;
  wire [31:0] T_1414_bits;
  wire [4:0] T_1414_rd;
  wire [4:0] T_1414_rs1;
  wire [4:0] T_1414_rs2;
  wire [4:0] T_1414_rs3;
  wire [4:0] T_1421;
  wire [4:0] T_1422;
  wire [31:0] T_1430_bits;
  wire [4:0] T_1430_rd;
  wire [4:0] T_1430_rs1;
  wire [4:0] T_1430_rs2;
  wire [4:0] T_1430_rs3;
  wire [31:0] T_1446_bits;
  wire [4:0] T_1446_rd;
  wire [4:0] T_1446_rs1;
  wire [4:0] T_1446_rs2;
  wire [4:0] T_1446_rs3;
  wire [31:0] T_1462_bits;
  wire [4:0] T_1462_rd;
  wire [4:0] T_1462_rs1;
  wire [4:0] T_1462_rs2;
  wire [4:0] T_1462_rs3;
  wire [31:0] T_1478_bits;
  wire [4:0] T_1478_rd;
  wire [4:0] T_1478_rs1;
  wire [4:0] T_1478_rs2;
  wire [4:0] T_1478_rs3;
  wire [31:0] T_1494_bits;
  wire [4:0] T_1494_rd;
  wire [4:0] T_1494_rs1;
  wire [4:0] T_1494_rs2;
  wire [4:0] T_1494_rs3;
  wire [31:0] T_1510_bits;
  wire [4:0] T_1510_rd;
  wire [4:0] T_1510_rs1;
  wire [4:0] T_1510_rs2;
  wire [4:0] T_1510_rs3;
  wire [31:0] T_1526_bits;
  wire [4:0] T_1526_rd;
  wire [4:0] T_1526_rs1;
  wire [4:0] T_1526_rs2;
  wire [4:0] T_1526_rs3;
  wire [31:0] T_1542_bits;
  wire [4:0] T_1542_rd;
  wire [4:0] T_1542_rs1;
  wire [4:0] T_1542_rs2;
  wire [4:0] T_1542_rs3;
  wire [2:0] T_1549;
  wire [4:0] T_1550;
  wire [4:0] T_1552;
  wire  T_1554;
  wire [4:0] T_1556;
  wire  T_1558;
  wire [4:0] T_1560;
  wire  T_1562;
  wire [4:0] T_1564;
  wire  T_1566;
  wire  T_1570;
  wire [31:0] T_1571_bits;
  wire [4:0] T_1571_rd;
  wire [4:0] T_1571_rs1;
  wire [4:0] T_1571_rs2;
  wire [4:0] T_1571_rs3;
  wire [31:0] T_1581_bits;
  wire [4:0] T_1581_rd;
  wire [4:0] T_1581_rs1;
  wire [4:0] T_1581_rs2;
  wire [4:0] T_1581_rs3;
  wire [31:0] T_1587_bits;
  wire [4:0] T_1587_rd;
  wire [4:0] T_1587_rs1;
  wire [4:0] T_1587_rs2;
  wire [4:0] T_1587_rs3;
  wire [31:0] T_1601_bits;
  wire [4:0] T_1601_rd;
  wire [4:0] T_1601_rs1;
  wire [4:0] T_1601_rs2;
  wire [4:0] T_1601_rs3;
  wire [31:0] T_1611_bits;
  wire [4:0] T_1611_rd;
  wire [4:0] T_1611_rs1;
  wire [4:0] T_1611_rs2;
  wire [4:0] T_1611_rs3;
  wire [31:0] T_1617_bits;
  wire [4:0] T_1617_rd;
  wire [4:0] T_1617_rs1;
  wire [4:0] T_1617_rs2;
  wire [4:0] T_1617_rs3;
  wire [31:0] T_1623_bits;
  wire [4:0] T_1623_rd;
  wire [4:0] T_1623_rs1;
  wire [4:0] T_1623_rs2;
  wire [4:0] T_1623_rs3;
  wire [31:0] T_1641_bits;
  wire [4:0] T_1641_rd;
  wire [4:0] T_1641_rs1;
  wire [4:0] T_1641_rs2;
  wire [4:0] T_1641_rs3;
  wire [31:0] T_1651_bits;
  wire [4:0] T_1651_rd;
  wire [4:0] T_1651_rs1;
  wire [4:0] T_1651_rs2;
  wire [4:0] T_1651_rs3;
  wire [31:0] T_1657_bits;
  wire [4:0] T_1657_rd;
  wire [4:0] T_1657_rs1;
  wire [4:0] T_1657_rs2;
  wire [4:0] T_1657_rs3;
  wire [31:0] T_1671_bits;
  wire [4:0] T_1671_rd;
  wire [4:0] T_1671_rs1;
  wire [4:0] T_1671_rs2;
  wire [4:0] T_1671_rs3;
  wire [31:0] T_1681_bits;
  wire [4:0] T_1681_rd;
  wire [4:0] T_1681_rs1;
  wire [4:0] T_1681_rs2;
  wire [4:0] T_1681_rs3;
  wire [31:0] T_1687_bits;
  wire [4:0] T_1687_rd;
  wire [4:0] T_1687_rs1;
  wire [4:0] T_1687_rs2;
  wire [4:0] T_1687_rs3;
  wire [31:0] T_1693_bits;
  wire [4:0] T_1693_rd;
  wire [4:0] T_1693_rs1;
  wire [4:0] T_1693_rs2;
  wire [4:0] T_1693_rs3;
  wire [31:0] T_1699_bits;
  wire [4:0] T_1699_rd;
  wire [4:0] T_1699_rs1;
  wire [4:0] T_1699_rs2;
  wire [4:0] T_1699_rs3;
  wire [31:0] T_1721_bits;
  wire [4:0] T_1721_rd;
  wire [4:0] T_1721_rs1;
  wire [4:0] T_1721_rs2;
  wire [4:0] T_1721_rs3;
  wire [31:0] T_1731_bits;
  wire [4:0] T_1731_rd;
  wire [4:0] T_1731_rs1;
  wire [4:0] T_1731_rs2;
  wire [4:0] T_1731_rs3;
  wire [31:0] T_1737_bits;
  wire [4:0] T_1737_rd;
  wire [4:0] T_1737_rs1;
  wire [4:0] T_1737_rs2;
  wire [4:0] T_1737_rs3;
  wire [31:0] T_1751_bits;
  wire [4:0] T_1751_rd;
  wire [4:0] T_1751_rs1;
  wire [4:0] T_1751_rs2;
  wire [4:0] T_1751_rs3;
  wire [31:0] T_1761_bits;
  wire [4:0] T_1761_rd;
  wire [4:0] T_1761_rs1;
  wire [4:0] T_1761_rs2;
  wire [4:0] T_1761_rs3;
  wire [31:0] T_1767_bits;
  wire [4:0] T_1767_rd;
  wire [4:0] T_1767_rs1;
  wire [4:0] T_1767_rs2;
  wire [4:0] T_1767_rs3;
  wire [31:0] T_1773_bits;
  wire [4:0] T_1773_rd;
  wire [4:0] T_1773_rs1;
  wire [4:0] T_1773_rs2;
  wire [4:0] T_1773_rs3;
  wire [31:0] T_1791_bits;
  wire [4:0] T_1791_rd;
  wire [4:0] T_1791_rs1;
  wire [4:0] T_1791_rs2;
  wire [4:0] T_1791_rs3;
  wire [31:0] T_1801_bits;
  wire [4:0] T_1801_rd;
  wire [4:0] T_1801_rs1;
  wire [4:0] T_1801_rs2;
  wire [4:0] T_1801_rs3;
  wire [31:0] T_1807_bits;
  wire [4:0] T_1807_rd;
  wire [4:0] T_1807_rs1;
  wire [4:0] T_1807_rs2;
  wire [4:0] T_1807_rs3;
  wire [31:0] T_1821_bits;
  wire [4:0] T_1821_rd;
  wire [4:0] T_1821_rs1;
  wire [4:0] T_1821_rs2;
  wire [4:0] T_1821_rs3;
  wire [31:0] T_1831_bits;
  wire [4:0] T_1831_rd;
  wire [4:0] T_1831_rs1;
  wire [4:0] T_1831_rs2;
  wire [4:0] T_1831_rs3;
  wire [31:0] T_1837_bits;
  wire [4:0] T_1837_rd;
  wire [4:0] T_1837_rs1;
  wire [4:0] T_1837_rs2;
  wire [4:0] T_1837_rs3;
  wire [31:0] T_1843_bits;
  wire [4:0] T_1843_rd;
  wire [4:0] T_1843_rs1;
  wire [4:0] T_1843_rs2;
  wire [4:0] T_1843_rs3;
  wire [31:0] T_1849_bits;
  wire [4:0] T_1849_rd;
  wire [4:0] T_1849_rs1;
  wire [4:0] T_1849_rs2;
  wire [4:0] T_1849_rs3;
  wire [31:0] T_1855_bits;
  wire [4:0] T_1855_rd;
  wire [4:0] T_1855_rs1;
  wire [4:0] T_1855_rs2;
  wire [4:0] T_1855_rs3;
  assign io_out_bits = T_1855_bits;
  assign io_out_rd = T_1855_rd;
  assign io_out_rs1 = T_1855_rs1;
  assign io_out_rs2 = T_1855_rs2;
  assign io_out_rs3 = T_1855_rs3;
  assign io_rvc = T_10;
  assign T_8 = io_in[1:0];
  assign T_10 = T_8 != 2'h3;
  assign T_11 = io_in[12:5];
  assign T_13 = T_11 != 8'h0;
  assign T_16 = T_13 ? 7'h13 : 7'h1f;
  assign T_17 = io_in[10:7];
  assign T_18 = io_in[12:11];
  assign T_19 = io_in[5];
  assign T_20 = io_in[6];
  assign T_22 = {T_20,2'h0};
  assign T_23 = {T_17,T_18};
  assign T_24 = {T_23,T_19};
  assign T_25 = {T_24,T_22};
  assign T_29 = io_in[4:2];
  assign T_30 = {2'h1,T_29};
  assign T_31 = {T_30,T_16};
  assign T_32 = {T_25,5'h2};
  assign T_33 = {T_32,3'h0};
  assign T_34 = {T_33,T_31};
  assign T_42 = io_in[31:27];
  assign T_49_bits = {{2'd0}, T_34};
  assign T_49_rd = T_30;
  assign T_49_rs1 = 5'h2;
  assign T_49_rs2 = T_30;
  assign T_49_rs3 = T_42;
  assign T_55 = io_in[6:5];
  assign T_56 = io_in[12:10];
  assign T_58 = {T_55,T_56};
  assign T_59 = {T_58,3'h0};
  assign T_61 = io_in[9:7];
  assign T_62 = {2'h1,T_61};
  assign T_68 = {T_30,7'h7};
  assign T_69 = {T_59,T_62};
  assign T_70 = {T_69,3'h3};
  assign T_71 = {T_70,T_68};
  assign T_88_bits = {{4'd0}, T_71};
  assign T_88_rd = T_30;
  assign T_88_rs1 = T_62;
  assign T_88_rs2 = T_30;
  assign T_88_rs3 = T_42;
  assign T_99 = {T_19,T_56};
  assign T_100 = {T_99,T_22};
  assign T_109 = {T_30,7'h3};
  assign T_110 = {T_100,T_62};
  assign T_111 = {T_110,3'h2};
  assign T_112 = {T_111,T_109};
  assign T_129_bits = {{5'd0}, T_112};
  assign T_129_rd = T_30;
  assign T_129_rs1 = T_62;
  assign T_129_rs2 = T_30;
  assign T_129_rs3 = T_42;
  assign T_151 = {T_70,T_109};
  assign T_168_bits = {{4'd0}, T_151};
  assign T_168_rd = T_30;
  assign T_168_rs1 = T_62;
  assign T_168_rs2 = T_30;
  assign T_168_rs3 = T_42;
  assign T_181 = T_100[6:5];
  assign T_196 = T_100[4:0];
  assign T_198 = {3'h2,T_196};
  assign T_199 = {T_198,7'h2f};
  assign T_200 = {T_181,T_30};
  assign T_201 = {T_200,T_62};
  assign T_202 = {T_201,T_199};
  assign T_219_bits = {{5'd0}, T_202};
  assign T_219_rd = T_30;
  assign T_219_rs1 = T_62;
  assign T_219_rs2 = T_30;
  assign T_219_rs3 = T_42;
  assign T_230 = T_59[7:5];
  assign T_243 = T_59[4:0];
  assign T_245 = {3'h3,T_243};
  assign T_246 = {T_245,7'h27};
  assign T_247 = {T_230,T_30};
  assign T_248 = {T_247,T_62};
  assign T_249 = {T_248,T_246};
  assign T_266_bits = {{4'd0}, T_249};
  assign T_266_rd = T_30;
  assign T_266_rs1 = T_62;
  assign T_266_rs2 = T_30;
  assign T_266_rs3 = T_42;
  assign T_297 = {T_198,7'h23};
  assign T_300 = {T_201,T_297};
  assign T_317_bits = {{5'd0}, T_300};
  assign T_317_rd = T_30;
  assign T_317_rs1 = T_62;
  assign T_317_rs2 = T_30;
  assign T_317_rs3 = T_42;
  assign T_344 = {T_245,7'h23};
  assign T_347 = {T_248,T_344};
  assign T_364_bits = {{4'd0}, T_347};
  assign T_364_rd = T_30;
  assign T_364_rs1 = T_62;
  assign T_364_rs2 = T_30;
  assign T_364_rs3 = T_42;
  assign T_370 = io_in[12];
  assign T_374 = T_370 ? 7'h7f : 7'h0;
  assign T_375 = io_in[6:2];
  assign T_376 = {T_374,T_375};
  assign T_377 = io_in[11:7];
  assign T_381 = {T_377,7'h13};
  assign T_382 = {T_376,T_377};
  assign T_383 = {T_382,3'h0};
  assign T_384 = {T_383,T_381};
  assign T_397_bits = T_384;
  assign T_397_rd = T_377;
  assign T_397_rs1 = T_377;
  assign T_397_rs2 = T_30;
  assign T_397_rs3 = T_42;
  assign T_405 = T_377 != 5'h0;
  assign T_408 = T_405 ? 7'h1b : 7'h1f;
  assign T_419 = {T_377,T_408};
  assign T_422 = {T_383,T_419};
  assign T_435_bits = T_422;
  assign T_435_rd = T_377;
  assign T_435_rs1 = T_377;
  assign T_435_rs2 = T_30;
  assign T_435_rs3 = T_42;
  assign T_453 = {T_376,5'h0};
  assign T_454 = {T_453,3'h0};
  assign T_455 = {T_454,T_381};
  assign T_468_bits = T_455;
  assign T_468_rd = T_377;
  assign T_468_rs1 = 5'h0;
  assign T_468_rs2 = T_30;
  assign T_468_rs3 = T_42;
  assign T_482 = T_376 != 12'h0;
  assign T_485 = T_482 ? 7'h37 : 7'h3f;
  assign T_490 = T_370 ? 15'h7fff : 15'h0;
  assign T_493 = {T_490,T_375};
  assign T_494 = {T_493,12'h0};
  assign T_495 = T_494[31:12];
  assign T_497 = {T_495,T_377};
  assign T_498 = {T_497,T_485};
  assign T_511_bits = T_498;
  assign T_511_rd = T_377;
  assign T_511_rs1 = T_377;
  assign T_511_rs2 = T_30;
  assign T_511_rs3 = T_42;
  assign T_519 = T_377 == 5'h0;
  assign T_522 = T_377 == 5'h2;
  assign T_523 = T_519 | T_522;
  assign T_535 = T_482 ? 7'h13 : 7'h1f;
  assign T_540 = T_370 ? 3'h7 : 3'h0;
  assign T_541 = io_in[4:3];
  assign T_543 = io_in[2];
  assign T_546 = {T_543,T_20};
  assign T_547 = {T_546,4'h0};
  assign T_548 = {T_540,T_541};
  assign T_549 = {T_548,T_19};
  assign T_550 = {T_549,T_547};
  assign T_554 = {T_377,T_535};
  assign T_555 = {T_550,T_377};
  assign T_556 = {T_555,3'h0};
  assign T_557 = {T_556,T_554};
  assign T_570_bits = T_557;
  assign T_570_rd = T_377;
  assign T_570_rs1 = T_377;
  assign T_570_rs2 = T_30;
  assign T_570_rs3 = T_42;
  assign T_576_bits = T_523 ? T_570_bits : T_511_bits;
  assign T_576_rd = T_523 ? T_570_rd : T_511_rd;
  assign T_576_rs1 = T_523 ? T_570_rs1 : T_511_rs1;
  assign T_576_rs2 = T_523 ? T_570_rs2 : T_511_rs2;
  assign T_576_rs3 = T_523 ? T_570_rs3 : T_511_rs3;
  assign T_584 = {T_370,T_375};
  assign T_593 = {T_62,7'h13};
  assign T_594 = {T_584,T_62};
  assign T_595 = {T_594,3'h5};
  assign T_596 = {T_595,T_593};
  assign GEN_0 = {{5'd0}, T_596};
  assign T_613 = GEN_0 | 31'h40000000;
  assign T_630 = {T_376,T_62};
  assign T_631 = {T_630,3'h7};
  assign T_632 = {T_631,T_593};
  assign T_643 = {T_370,T_55};
  assign T_645 = T_643 & 3'h3;
  assign T_647 = T_643 >= 3'h4;
  assign T_649 = T_645 & 3'h1;
  assign T_651 = T_645 >= 3'h2;
  assign T_655 = T_649 >= 3'h1;
  assign T_656 = T_655 ? 2'h3 : 2'h2;
  assign T_662 = T_651 ? T_656 : 2'h0;
  assign T_671 = T_655 ? 3'h7 : 3'h6;
  assign T_676 = T_655 ? 3'h4 : 3'h0;
  assign T_677 = T_651 ? T_671 : T_676;
  assign T_678 = T_647 ? {{1'd0}, T_662} : T_677;
  assign T_681 = T_55 == 2'h0;
  assign T_684 = T_681 ? 31'h40000000 : 31'h0;
  assign T_688 = T_370 ? 7'h3b : 7'h33;
  assign T_698 = {T_62,T_688};
  assign T_699 = {T_30,T_62};
  assign T_700 = {T_699,T_678};
  assign T_701 = {T_700,T_698};
  assign GEN_1 = {{6'd0}, T_701};
  assign T_702 = GEN_1 | T_684;
  assign T_703 = io_in[11:10];
  assign T_705 = T_703 & 2'h1;
  assign T_707 = T_703 >= 2'h2;
  assign T_711 = T_705 >= 2'h1;
  assign T_712 = T_711 ? {{1'd0}, T_702} : T_632;
  assign T_717 = T_711 ? T_613 : {{5'd0}, T_596};
  assign T_718 = T_707 ? T_712 : {{1'd0}, T_717};
  assign T_735_bits = T_718;
  assign T_735_rd = T_62;
  assign T_735_rs1 = T_62;
  assign T_735_rs2 = T_30;
  assign T_735_rs3 = T_42;
  assign T_745 = T_370 ? 10'h3ff : 10'h0;
  assign T_746 = io_in[8];
  assign T_747 = io_in[10:9];
  assign T_749 = io_in[7];
  assign T_751 = io_in[11];
  assign T_752 = io_in[5:3];
  assign T_754 = {T_752,1'h0};
  assign T_755 = {T_543,T_751};
  assign T_756 = {T_755,T_754};
  assign T_757 = {T_20,T_749};
  assign T_758 = {T_745,T_746};
  assign T_759 = {T_758,T_747};
  assign T_760 = {T_759,T_757};
  assign T_761 = {T_760,T_756};
  assign T_762 = T_761[20];
  assign T_784 = T_761[10:1];
  assign T_806 = T_761[11];
  assign T_828 = T_761[19:12];
  assign T_831 = {T_828,5'h0};
  assign T_832 = {T_831,7'h6f};
  assign T_833 = {T_762,T_784};
  assign T_834 = {T_833,T_806};
  assign T_835 = {T_834,T_832};
  assign T_850_bits = T_835;
  assign T_850_rd = 5'h0;
  assign T_850_rs1 = T_62;
  assign T_850_rs2 = T_30;
  assign T_850_rs3 = T_42;
  assign T_860 = T_370 ? 5'h1f : 5'h0;
  assign T_866 = {T_703,T_541};
  assign T_867 = {T_866,1'h0};
  assign T_868 = {T_860,T_55};
  assign T_869 = {T_868,T_543};
  assign T_870 = {T_869,T_867};
  assign T_871 = T_870[12];
  assign T_887 = T_870[10:5];
  assign T_908 = T_870[4:1];
  assign T_924 = T_870[11];
  assign T_926 = {T_924,7'h63};
  assign T_927 = {3'h0,T_908};
  assign T_928 = {T_927,T_926};
  assign T_929 = {5'h0,T_62};
  assign T_930 = {T_871,T_887};
  assign T_931 = {T_930,T_929};
  assign T_932 = {T_931,T_928};
  assign T_947_bits = T_932;
  assign T_947_rd = T_62;
  assign T_947_rs1 = T_62;
  assign T_947_rs2 = 5'h0;
  assign T_947_rs3 = T_42;
  assign T_1024 = {3'h1,T_908};
  assign T_1025 = {T_1024,T_926};
  assign T_1029 = {T_931,T_1025};
  assign T_1042_bits = T_1029;
  assign T_1042_rd = 5'h0;
  assign T_1042_rs1 = T_62;
  assign T_1042_rs2 = 5'h0;
  assign T_1042_rs3 = T_42;
  assign T_1056 = {T_584,T_377};
  assign T_1057 = {T_1056,3'h1};
  assign T_1058 = {T_1057,T_381};
  assign T_1069_bits = {{6'd0}, T_1058};
  assign T_1069_rd = T_377;
  assign T_1069_rs1 = T_377;
  assign T_1069_rs2 = T_375;
  assign T_1069_rs3 = T_42;
  assign T_1079 = {T_55,3'h0};
  assign T_1080 = {T_29,T_370};
  assign T_1081 = {T_1080,T_1079};
  assign T_1086 = {T_377,7'h7};
  assign T_1087 = {T_1081,5'h2};
  assign T_1088 = {T_1087,3'h3};
  assign T_1089 = {T_1088,T_1086};
  assign T_1100_bits = {{3'd0}, T_1089};
  assign T_1100_rd = T_377;
  assign T_1100_rs1 = 5'h2;
  assign T_1100_rs2 = T_375;
  assign T_1100_rs3 = T_42;
  assign T_1106 = io_in[3:2];
  assign T_1108 = io_in[6:4];
  assign T_1110 = {T_1108,2'h0};
  assign T_1111 = {T_1106,T_370};
  assign T_1112 = {T_1111,T_1110};
  assign T_1117 = {T_377,7'h3};
  assign T_1118 = {T_1112,5'h2};
  assign T_1119 = {T_1118,3'h2};
  assign T_1120 = {T_1119,T_1117};
  assign T_1131_bits = {{4'd0}, T_1120};
  assign T_1131_rd = T_377;
  assign T_1131_rs1 = 5'h2;
  assign T_1131_rs2 = T_375;
  assign T_1131_rs3 = T_42;
  assign T_1151 = {T_1088,T_1117};
  assign T_1162_bits = {{3'd0}, T_1151};
  assign T_1162_rd = T_377;
  assign T_1162_rs1 = 5'h2;
  assign T_1162_rs2 = T_375;
  assign T_1162_rs3 = T_42;
  assign T_1173 = {T_377,7'h33};
  assign T_1174 = {T_375,5'h0};
  assign T_1175 = {T_1174,3'h0};
  assign T_1176 = {T_1175,T_1173};
  assign T_1187_bits = {{7'd0}, T_1176};
  assign T_1187_rd = T_377;
  assign T_1187_rs1 = 5'h0;
  assign T_1187_rs2 = T_375;
  assign T_1187_rs3 = T_42;
  assign T_1199 = {T_375,T_377};
  assign T_1200 = {T_1199,3'h0};
  assign T_1201 = {T_1200,T_1173};
  assign T_1212_bits = {{7'd0}, T_1201};
  assign T_1212_rd = T_377;
  assign T_1212_rs1 = T_377;
  assign T_1212_rs2 = T_375;
  assign T_1212_rs3 = T_42;
  assign T_1226 = {T_1200,12'h67};
  assign T_1227 = T_1226[24:7];
  assign T_1229 = {T_1227,7'h1f};
  assign T_1233 = T_405 ? T_1226 : T_1229;
  assign T_1244_bits = {{7'd0}, T_1233};
  assign T_1244_rd = 5'h0;
  assign T_1244_rs1 = T_377;
  assign T_1244_rs2 = T_375;
  assign T_1244_rs3 = T_42;
  assign T_1252 = T_375 != 5'h0;
  assign T_1253_bits = T_1252 ? T_1187_bits : T_1244_bits;
  assign T_1253_rd = T_1252 ? T_1187_rd : T_1244_rd;
  assign T_1253_rs1 = T_1252 ? T_1187_rs1 : T_1244_rs1;
  assign T_1253_rs2 = T_1252 ? T_1187_rs2 : T_1244_rs2;
  assign T_1253_rs3 = T_1252 ? T_1187_rs3 : T_1244_rs3;
  assign T_1267 = {T_1200,12'he7};
  assign T_1270 = {T_1227,7'h73};
  assign T_1272 = T_1270 | 25'h100000;
  assign T_1276 = T_405 ? T_1267 : T_1272;
  assign T_1287_bits = {{7'd0}, T_1276};
  assign T_1287_rd = 5'h1;
  assign T_1287_rs1 = T_377;
  assign T_1287_rs2 = T_375;
  assign T_1287_rs3 = T_42;
  assign T_1296_bits = T_1252 ? T_1212_bits : T_1287_bits;
  assign T_1296_rd = T_1252 ? T_1212_rd : T_1287_rd;
  assign T_1296_rs1 = T_1252 ? T_1212_rs1 : T_1287_rs1;
  assign T_1296_rs2 = T_1252 ? T_1212_rs2 : T_1287_rs2;
  assign T_1296_rs3 = T_1252 ? T_1212_rs3 : T_1287_rs3;
  assign T_1303_bits = T_370 ? T_1296_bits : T_1253_bits;
  assign T_1303_rd = T_370 ? T_1296_rd : T_1253_rd;
  assign T_1303_rs1 = T_370 ? T_1296_rs1 : T_1253_rs1;
  assign T_1303_rs2 = T_370 ? T_1296_rs2 : T_1253_rs2;
  assign T_1303_rs3 = T_370 ? T_1296_rs3 : T_1253_rs3;
  assign T_1312 = {T_61,T_56};
  assign T_1313 = {T_1312,3'h0};
  assign T_1314 = T_1313[8:5];
  assign T_1323 = T_1313[4:0];
  assign T_1325 = {3'h3,T_1323};
  assign T_1326 = {T_1325,7'h27};
  assign T_1327 = {T_1314,T_375};
  assign T_1328 = {T_1327,5'h2};
  assign T_1329 = {T_1328,T_1326};
  assign T_1340_bits = {{3'd0}, T_1329};
  assign T_1340_rd = T_377;
  assign T_1340_rs1 = 5'h2;
  assign T_1340_rs2 = T_375;
  assign T_1340_rs3 = T_42;
  assign T_1346 = io_in[8:7];
  assign T_1347 = io_in[12:9];
  assign T_1349 = {T_1346,T_1347};
  assign T_1350 = {T_1349,2'h0};
  assign T_1351 = T_1350[7:5];
  assign T_1360 = T_1350[4:0];
  assign T_1362 = {3'h2,T_1360};
  assign T_1363 = {T_1362,7'h23};
  assign T_1364 = {T_1351,T_375};
  assign T_1365 = {T_1364,5'h2};
  assign T_1366 = {T_1365,T_1363};
  assign T_1377_bits = {{4'd0}, T_1366};
  assign T_1377_rd = T_377;
  assign T_1377_rs1 = 5'h2;
  assign T_1377_rs2 = T_375;
  assign T_1377_rs3 = T_42;
  assign T_1400 = {T_1325,7'h23};
  assign T_1403 = {T_1328,T_1400};
  assign T_1414_bits = {{3'd0}, T_1403};
  assign T_1414_rd = T_377;
  assign T_1414_rs1 = 5'h2;
  assign T_1414_rs2 = T_375;
  assign T_1414_rs3 = T_42;
  assign T_1421 = io_in[19:15];
  assign T_1422 = io_in[24:20];
  assign T_1430_bits = io_in;
  assign T_1430_rd = T_377;
  assign T_1430_rs1 = T_1421;
  assign T_1430_rs2 = T_1422;
  assign T_1430_rs3 = T_42;
  assign T_1446_bits = io_in;
  assign T_1446_rd = T_377;
  assign T_1446_rs1 = T_1421;
  assign T_1446_rs2 = T_1422;
  assign T_1446_rs3 = T_42;
  assign T_1462_bits = io_in;
  assign T_1462_rd = T_377;
  assign T_1462_rs1 = T_1421;
  assign T_1462_rs2 = T_1422;
  assign T_1462_rs3 = T_42;
  assign T_1478_bits = io_in;
  assign T_1478_rd = T_377;
  assign T_1478_rs1 = T_1421;
  assign T_1478_rs2 = T_1422;
  assign T_1478_rs3 = T_42;
  assign T_1494_bits = io_in;
  assign T_1494_rd = T_377;
  assign T_1494_rs1 = T_1421;
  assign T_1494_rs2 = T_1422;
  assign T_1494_rs3 = T_42;
  assign T_1510_bits = io_in;
  assign T_1510_rd = T_377;
  assign T_1510_rs1 = T_1421;
  assign T_1510_rs2 = T_1422;
  assign T_1510_rs3 = T_42;
  assign T_1526_bits = io_in;
  assign T_1526_rd = T_377;
  assign T_1526_rs1 = T_1421;
  assign T_1526_rs2 = T_1422;
  assign T_1526_rs3 = T_42;
  assign T_1542_bits = io_in;
  assign T_1542_rd = T_377;
  assign T_1542_rs1 = T_1421;
  assign T_1542_rs2 = T_1422;
  assign T_1542_rs3 = T_42;
  assign T_1549 = io_in[15:13];
  assign T_1550 = {T_8,T_1549};
  assign T_1552 = T_1550 & 5'hf;
  assign T_1554 = T_1550 >= 5'h10;
  assign T_1556 = T_1552 & 5'h7;
  assign T_1558 = T_1552 >= 5'h8;
  assign T_1560 = T_1556 & 5'h3;
  assign T_1562 = T_1556 >= 5'h4;
  assign T_1564 = T_1560 & 5'h1;
  assign T_1566 = T_1560 >= 5'h2;
  assign T_1570 = T_1564 >= 5'h1;
  assign T_1571_bits = T_1570 ? T_1542_bits : T_1526_bits;
  assign T_1571_rd = T_1570 ? T_1542_rd : T_1526_rd;
  assign T_1571_rs1 = T_1570 ? T_1542_rs1 : T_1526_rs1;
  assign T_1571_rs2 = T_1570 ? T_1542_rs2 : T_1526_rs2;
  assign T_1571_rs3 = T_1570 ? T_1542_rs3 : T_1526_rs3;
  assign T_1581_bits = T_1570 ? T_1510_bits : T_1494_bits;
  assign T_1581_rd = T_1570 ? T_1510_rd : T_1494_rd;
  assign T_1581_rs1 = T_1570 ? T_1510_rs1 : T_1494_rs1;
  assign T_1581_rs2 = T_1570 ? T_1510_rs2 : T_1494_rs2;
  assign T_1581_rs3 = T_1570 ? T_1510_rs3 : T_1494_rs3;
  assign T_1587_bits = T_1566 ? T_1571_bits : T_1581_bits;
  assign T_1587_rd = T_1566 ? T_1571_rd : T_1581_rd;
  assign T_1587_rs1 = T_1566 ? T_1571_rs1 : T_1581_rs1;
  assign T_1587_rs2 = T_1566 ? T_1571_rs2 : T_1581_rs2;
  assign T_1587_rs3 = T_1566 ? T_1571_rs3 : T_1581_rs3;
  assign T_1601_bits = T_1570 ? T_1478_bits : T_1462_bits;
  assign T_1601_rd = T_1570 ? T_1478_rd : T_1462_rd;
  assign T_1601_rs1 = T_1570 ? T_1478_rs1 : T_1462_rs1;
  assign T_1601_rs2 = T_1570 ? T_1478_rs2 : T_1462_rs2;
  assign T_1601_rs3 = T_1570 ? T_1478_rs3 : T_1462_rs3;
  assign T_1611_bits = T_1570 ? T_1446_bits : T_1430_bits;
  assign T_1611_rd = T_1570 ? T_1446_rd : T_1430_rd;
  assign T_1611_rs1 = T_1570 ? T_1446_rs1 : T_1430_rs1;
  assign T_1611_rs2 = T_1570 ? T_1446_rs2 : T_1430_rs2;
  assign T_1611_rs3 = T_1570 ? T_1446_rs3 : T_1430_rs3;
  assign T_1617_bits = T_1566 ? T_1601_bits : T_1611_bits;
  assign T_1617_rd = T_1566 ? T_1601_rd : T_1611_rd;
  assign T_1617_rs1 = T_1566 ? T_1601_rs1 : T_1611_rs1;
  assign T_1617_rs2 = T_1566 ? T_1601_rs2 : T_1611_rs2;
  assign T_1617_rs3 = T_1566 ? T_1601_rs3 : T_1611_rs3;
  assign T_1623_bits = T_1562 ? T_1587_bits : T_1617_bits;
  assign T_1623_rd = T_1562 ? T_1587_rd : T_1617_rd;
  assign T_1623_rs1 = T_1562 ? T_1587_rs1 : T_1617_rs1;
  assign T_1623_rs2 = T_1562 ? T_1587_rs2 : T_1617_rs2;
  assign T_1623_rs3 = T_1562 ? T_1587_rs3 : T_1617_rs3;
  assign T_1641_bits = T_1570 ? T_1414_bits : T_1377_bits;
  assign T_1641_rd = T_1570 ? T_1414_rd : T_1377_rd;
  assign T_1641_rs1 = T_1570 ? T_1414_rs1 : T_1377_rs1;
  assign T_1641_rs2 = T_1570 ? T_1414_rs2 : T_1377_rs2;
  assign T_1641_rs3 = T_1570 ? T_1414_rs3 : T_1377_rs3;
  assign T_1651_bits = T_1570 ? T_1340_bits : T_1303_bits;
  assign T_1651_rd = T_1570 ? T_1340_rd : T_1303_rd;
  assign T_1651_rs1 = T_1570 ? T_1340_rs1 : T_1303_rs1;
  assign T_1651_rs2 = T_1570 ? T_1340_rs2 : T_1303_rs2;
  assign T_1651_rs3 = T_1570 ? T_1340_rs3 : T_1303_rs3;
  assign T_1657_bits = T_1566 ? T_1641_bits : T_1651_bits;
  assign T_1657_rd = T_1566 ? T_1641_rd : T_1651_rd;
  assign T_1657_rs1 = T_1566 ? T_1641_rs1 : T_1651_rs1;
  assign T_1657_rs2 = T_1566 ? T_1641_rs2 : T_1651_rs2;
  assign T_1657_rs3 = T_1566 ? T_1641_rs3 : T_1651_rs3;
  assign T_1671_bits = T_1570 ? T_1162_bits : T_1131_bits;
  assign T_1671_rd = T_1570 ? T_1162_rd : T_1131_rd;
  assign T_1671_rs1 = T_1570 ? T_1162_rs1 : T_1131_rs1;
  assign T_1671_rs2 = T_1570 ? T_1162_rs2 : T_1131_rs2;
  assign T_1671_rs3 = T_1570 ? T_1162_rs3 : T_1131_rs3;
  assign T_1681_bits = T_1570 ? T_1100_bits : T_1069_bits;
  assign T_1681_rd = T_1570 ? T_1100_rd : T_1069_rd;
  assign T_1681_rs1 = T_1570 ? T_1100_rs1 : T_1069_rs1;
  assign T_1681_rs2 = T_1570 ? T_1100_rs2 : T_1069_rs2;
  assign T_1681_rs3 = T_1570 ? T_1100_rs3 : T_1069_rs3;
  assign T_1687_bits = T_1566 ? T_1671_bits : T_1681_bits;
  assign T_1687_rd = T_1566 ? T_1671_rd : T_1681_rd;
  assign T_1687_rs1 = T_1566 ? T_1671_rs1 : T_1681_rs1;
  assign T_1687_rs2 = T_1566 ? T_1671_rs2 : T_1681_rs2;
  assign T_1687_rs3 = T_1566 ? T_1671_rs3 : T_1681_rs3;
  assign T_1693_bits = T_1562 ? T_1657_bits : T_1687_bits;
  assign T_1693_rd = T_1562 ? T_1657_rd : T_1687_rd;
  assign T_1693_rs1 = T_1562 ? T_1657_rs1 : T_1687_rs1;
  assign T_1693_rs2 = T_1562 ? T_1657_rs2 : T_1687_rs2;
  assign T_1693_rs3 = T_1562 ? T_1657_rs3 : T_1687_rs3;
  assign T_1699_bits = T_1558 ? T_1623_bits : T_1693_bits;
  assign T_1699_rd = T_1558 ? T_1623_rd : T_1693_rd;
  assign T_1699_rs1 = T_1558 ? T_1623_rs1 : T_1693_rs1;
  assign T_1699_rs2 = T_1558 ? T_1623_rs2 : T_1693_rs2;
  assign T_1699_rs3 = T_1558 ? T_1623_rs3 : T_1693_rs3;
  assign T_1721_bits = T_1570 ? T_1042_bits : T_947_bits;
  assign T_1721_rd = T_1570 ? T_1042_rd : T_947_rd;
  assign T_1721_rs1 = T_1570 ? T_1042_rs1 : T_947_rs1;
  assign T_1721_rs2 = T_1570 ? T_1042_rs2 : T_947_rs2;
  assign T_1721_rs3 = T_1570 ? T_1042_rs3 : T_947_rs3;
  assign T_1731_bits = T_1570 ? T_850_bits : T_735_bits;
  assign T_1731_rd = T_1570 ? T_850_rd : T_735_rd;
  assign T_1731_rs1 = T_1570 ? T_850_rs1 : T_735_rs1;
  assign T_1731_rs2 = T_1570 ? T_850_rs2 : T_735_rs2;
  assign T_1731_rs3 = T_1570 ? T_850_rs3 : T_735_rs3;
  assign T_1737_bits = T_1566 ? T_1721_bits : T_1731_bits;
  assign T_1737_rd = T_1566 ? T_1721_rd : T_1731_rd;
  assign T_1737_rs1 = T_1566 ? T_1721_rs1 : T_1731_rs1;
  assign T_1737_rs2 = T_1566 ? T_1721_rs2 : T_1731_rs2;
  assign T_1737_rs3 = T_1566 ? T_1721_rs3 : T_1731_rs3;
  assign T_1751_bits = T_1570 ? T_576_bits : T_468_bits;
  assign T_1751_rd = T_1570 ? T_576_rd : T_468_rd;
  assign T_1751_rs1 = T_1570 ? T_576_rs1 : T_468_rs1;
  assign T_1751_rs2 = T_1570 ? T_576_rs2 : T_468_rs2;
  assign T_1751_rs3 = T_1570 ? T_576_rs3 : T_468_rs3;
  assign T_1761_bits = T_1570 ? T_435_bits : T_397_bits;
  assign T_1761_rd = T_1570 ? T_435_rd : T_397_rd;
  assign T_1761_rs1 = T_1570 ? T_435_rs1 : T_397_rs1;
  assign T_1761_rs2 = T_1570 ? T_435_rs2 : T_397_rs2;
  assign T_1761_rs3 = T_1570 ? T_435_rs3 : T_397_rs3;
  assign T_1767_bits = T_1566 ? T_1751_bits : T_1761_bits;
  assign T_1767_rd = T_1566 ? T_1751_rd : T_1761_rd;
  assign T_1767_rs1 = T_1566 ? T_1751_rs1 : T_1761_rs1;
  assign T_1767_rs2 = T_1566 ? T_1751_rs2 : T_1761_rs2;
  assign T_1767_rs3 = T_1566 ? T_1751_rs3 : T_1761_rs3;
  assign T_1773_bits = T_1562 ? T_1737_bits : T_1767_bits;
  assign T_1773_rd = T_1562 ? T_1737_rd : T_1767_rd;
  assign T_1773_rs1 = T_1562 ? T_1737_rs1 : T_1767_rs1;
  assign T_1773_rs2 = T_1562 ? T_1737_rs2 : T_1767_rs2;
  assign T_1773_rs3 = T_1562 ? T_1737_rs3 : T_1767_rs3;
  assign T_1791_bits = T_1570 ? T_364_bits : T_317_bits;
  assign T_1791_rd = T_1570 ? T_364_rd : T_317_rd;
  assign T_1791_rs1 = T_1570 ? T_364_rs1 : T_317_rs1;
  assign T_1791_rs2 = T_1570 ? T_364_rs2 : T_317_rs2;
  assign T_1791_rs3 = T_1570 ? T_364_rs3 : T_317_rs3;
  assign T_1801_bits = T_1570 ? T_266_bits : T_219_bits;
  assign T_1801_rd = T_1570 ? T_266_rd : T_219_rd;
  assign T_1801_rs1 = T_1570 ? T_266_rs1 : T_219_rs1;
  assign T_1801_rs2 = T_1570 ? T_266_rs2 : T_219_rs2;
  assign T_1801_rs3 = T_1570 ? T_266_rs3 : T_219_rs3;
  assign T_1807_bits = T_1566 ? T_1791_bits : T_1801_bits;
  assign T_1807_rd = T_1566 ? T_1791_rd : T_1801_rd;
  assign T_1807_rs1 = T_1566 ? T_1791_rs1 : T_1801_rs1;
  assign T_1807_rs2 = T_1566 ? T_1791_rs2 : T_1801_rs2;
  assign T_1807_rs3 = T_1566 ? T_1791_rs3 : T_1801_rs3;
  assign T_1821_bits = T_1570 ? T_168_bits : T_129_bits;
  assign T_1821_rd = T_1570 ? T_168_rd : T_129_rd;
  assign T_1821_rs1 = T_1570 ? T_168_rs1 : T_129_rs1;
  assign T_1821_rs2 = T_1570 ? T_168_rs2 : T_129_rs2;
  assign T_1821_rs3 = T_1570 ? T_168_rs3 : T_129_rs3;
  assign T_1831_bits = T_1570 ? T_88_bits : T_49_bits;
  assign T_1831_rd = T_1570 ? T_88_rd : T_49_rd;
  assign T_1831_rs1 = T_1570 ? T_88_rs1 : T_49_rs1;
  assign T_1831_rs2 = T_1570 ? T_88_rs2 : T_49_rs2;
  assign T_1831_rs3 = T_1570 ? T_88_rs3 : T_49_rs3;
  assign T_1837_bits = T_1566 ? T_1821_bits : T_1831_bits;
  assign T_1837_rd = T_1566 ? T_1821_rd : T_1831_rd;
  assign T_1837_rs1 = T_1566 ? T_1821_rs1 : T_1831_rs1;
  assign T_1837_rs2 = T_1566 ? T_1821_rs2 : T_1831_rs2;
  assign T_1837_rs3 = T_1566 ? T_1821_rs3 : T_1831_rs3;
  assign T_1843_bits = T_1562 ? T_1807_bits : T_1837_bits;
  assign T_1843_rd = T_1562 ? T_1807_rd : T_1837_rd;
  assign T_1843_rs1 = T_1562 ? T_1807_rs1 : T_1837_rs1;
  assign T_1843_rs2 = T_1562 ? T_1807_rs2 : T_1837_rs2;
  assign T_1843_rs3 = T_1562 ? T_1807_rs3 : T_1837_rs3;
  assign T_1849_bits = T_1558 ? T_1773_bits : T_1843_bits;
  assign T_1849_rd = T_1558 ? T_1773_rd : T_1843_rd;
  assign T_1849_rs1 = T_1558 ? T_1773_rs1 : T_1843_rs1;
  assign T_1849_rs2 = T_1558 ? T_1773_rs2 : T_1843_rs2;
  assign T_1849_rs3 = T_1558 ? T_1773_rs3 : T_1843_rs3;
  assign T_1855_bits = T_1554 ? T_1699_bits : T_1849_bits;
  assign T_1855_rd = T_1554 ? T_1699_rd : T_1849_rd;
  assign T_1855_rs1 = T_1554 ? T_1699_rs1 : T_1849_rs1;
  assign T_1855_rs2 = T_1554 ? T_1699_rs2 : T_1849_rs2;
  assign T_1855_rs3 = T_1554 ? T_1699_rs3 : T_1849_rs3;
endmodule
module IBuf(
  input   clk,
  input   reset,
  output  io_imem_ready,
  input   io_imem_valid,
  input   io_imem_bits_btb_valid,
  input   io_imem_bits_btb_bits_taken,
  input  [1:0] io_imem_bits_btb_bits_mask,
  input   io_imem_bits_btb_bits_bridx,
  input  [38:0] io_imem_bits_btb_bits_target,
  input   io_imem_bits_btb_bits_entry,
  input   io_imem_bits_btb_bits_bht_history,
  input  [1:0] io_imem_bits_btb_bits_bht_value,
  input  [39:0] io_imem_bits_pc,
  input  [31:0] io_imem_bits_data,
  input  [1:0] io_imem_bits_mask,
  input   io_imem_bits_xcpt_if,
  input   io_imem_bits_replay,
  input   io_kill,
  output [39:0] io_pc,
  output  io_btb_resp_taken,
  output [1:0] io_btb_resp_mask,
  output  io_btb_resp_bridx,
  output [38:0] io_btb_resp_target,
  output  io_btb_resp_entry,
  output  io_btb_resp_bht_history,
  output [1:0] io_btb_resp_bht_value,
  input   io_inst_0_ready,
  output  io_inst_0_valid,
  output  io_inst_0_bits_pf0,
  output  io_inst_0_bits_pf1,
  output  io_inst_0_bits_replay,
  output  io_inst_0_bits_btb_hit,
  output  io_inst_0_bits_rvc,
  output [31:0] io_inst_0_bits_inst_bits,
  output [4:0] io_inst_0_bits_inst_rd,
  output [4:0] io_inst_0_bits_inst_rs1,
  output [4:0] io_inst_0_bits_inst_rs2,
  output [4:0] io_inst_0_bits_inst_rs3
);
  reg  nBufValid;
  reg [31:0] GEN_33;
  reg  buf_btb_valid;
  reg [31:0] GEN_34;
  reg  buf_btb_bits_taken;
  reg [31:0] GEN_35;
  reg [1:0] buf_btb_bits_mask;
  reg [31:0] GEN_36;
  reg  buf_btb_bits_bridx;
  reg [31:0] GEN_37;
  reg [38:0] buf_btb_bits_target;
  reg [63:0] GEN_38;
  reg  buf_btb_bits_entry;
  reg [31:0] GEN_43;
  reg  buf_btb_bits_bht_history;
  reg [31:0] GEN_44;
  reg [1:0] buf_btb_bits_bht_value;
  reg [31:0] GEN_48;
  reg [39:0] buf_pc;
  reg [63:0] GEN_51;
  reg [31:0] buf_data;
  reg [31:0] GEN_52;
  reg [1:0] buf_mask;
  reg [31:0] GEN_53;
  reg  buf_xcpt_if;
  reg [31:0] GEN_54;
  reg  buf_replay;
  reg [31:0] GEN_55;
  reg  ibufBTBHit;
  reg [31:0] GEN_56;
  reg  ibufBTBResp_taken;
  reg [31:0] GEN_57;
  reg [1:0] ibufBTBResp_mask;
  reg [31:0] GEN_58;
  reg  ibufBTBResp_bridx;
  reg [31:0] GEN_59;
  reg [38:0] ibufBTBResp_target;
  reg [63:0] GEN_60;
  reg  ibufBTBResp_entry;
  reg [31:0] GEN_61;
  reg  ibufBTBResp_bht_history;
  reg [31:0] GEN_62;
  reg [1:0] ibufBTBResp_bht_value;
  reg [31:0] GEN_63;
  wire  pcWordBits;
  wire [1:0] nReady;
  wire  T_375;
  wire [1:0] T_377;
  wire [1:0] T_379;
  wire [1:0] GEN_31;
  wire [2:0] T_380;
  wire [1:0] nIC;
  wire [1:0] GEN_32;
  wire [2:0] T_381;
  wire [1:0] nICReady;
  wire [1:0] T_383;
  wire [2:0] T_384;
  wire [1:0] nValid;
  wire  T_385;
  wire  T_386;
  wire [2:0] T_388;
  wire [1:0] T_389;
  wire  T_390;
  wire  T_391;
  wire  T_392;
  wire [2:0] T_395;
  wire [1:0] T_396;
  wire [1:0] T_397;
  wire  T_399;
  wire  T_400;
  wire  T_401;
  wire  T_406;
  wire [2:0] T_407;
  wire [1:0] T_408;
  wire [15:0] T_411;
  wire [31:0] T_412;
  wire [63:0] T_413;
  wire [5:0] GEN_39;
  wire [5:0] T_414;
  wire [63:0] T_415;
  wire [15:0] T_416;
  wire [39:0] T_418;
  wire [2:0] GEN_40;
  wire [2:0] T_419;
  wire [39:0] GEN_41;
  wire [40:0] T_420;
  wire [39:0] T_421;
  wire [39:0] T_422;
  wire [39:0] T_423;
  wire [1:0] GEN_42;
  wire [2:0] T_424;
  wire [1:0] T_425;
  wire  GEN_0;
  wire [1:0] GEN_1;
  wire [1:0] GEN_2;
  wire [38:0] GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire [1:0] GEN_6;
  wire [1:0] GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire [1:0] GEN_10;
  wire  GEN_11;
  wire [38:0] GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [1:0] GEN_15;
  wire [39:0] GEN_16;
  wire [31:0] GEN_17;
  wire [1:0] GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [38:0] GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire [1:0] GEN_28;
  wire [1:0] GEN_29;
  wire [2:0] T_428;
  wire [1:0] T_429;
  wire [2:0] T_430;
  wire [1:0] T_431;
  wire [15:0] T_432;
  wire [31:0] T_433;
  wire [63:0] T_434;
  wire [15:0] T_435;
  wire [31:0] T_436;
  wire [63:0] T_437;
  wire [127:0] T_438;
  wire [5:0] GEN_45;
  wire [5:0] T_439;
  wire [190:0] GEN_46;
  wire [190:0] T_440;
  wire [31:0] icData;
  wire [4:0] GEN_47;
  wire [4:0] T_443;
  wire [62:0] T_444;
  wire [31:0] icMask;
  wire [31:0] T_445;
  wire [31:0] T_446;
  wire [31:0] T_447;
  wire [31:0] inst;
  wire [3:0] T_449;
  wire [4:0] T_451;
  wire [3:0] T_452;
  wire [1:0] valid;
  wire [1:0] T_454;
  wire [2:0] T_456;
  wire [1:0] bufMask;
  wire [1:0] T_458;
  wire [1:0] T_459;
  wire [1:0] T_461;
  wire [1:0] T_462;
  wire [1:0] xcpt_if;
  wire [1:0] T_464;
  wire [1:0] T_467;
  wire [1:0] T_468;
  wire [1:0] ic_replay;
  wire [1:0] T_470;
  wire [1:0] ibufBTBHitMask;
  wire [1:0] T_472;
  wire [2:0] T_473;
  wire [1:0] T_474;
  wire [3:0] T_476;
  wire [3:0] icBTBHitMask;
  wire [1:0] T_478;
  wire [3:0] GEN_49;
  wire [3:0] T_480;
  wire [3:0] GEN_50;
  wire [3:0] btbHitMask;
  wire  T_483;
  wire  T_484_taken;
  wire [1:0] T_484_mask;
  wire  T_484_bridx;
  wire [38:0] T_484_target;
  wire  T_484_entry;
  wire  T_484_bht_history;
  wire [1:0] T_484_bht_value;
  wire  T_494;
  wire [39:0] T_495;
  wire  RVCExpander_1_clk;
  wire  RVCExpander_1_reset;
  wire [31:0] RVCExpander_1_io_in;
  wire [31:0] RVCExpander_1_io_out_bits;
  wire [4:0] RVCExpander_1_io_out_rd;
  wire [4:0] RVCExpander_1_io_out_rs1;
  wire [4:0] RVCExpander_1_io_out_rs2;
  wire [4:0] RVCExpander_1_io_out_rs3;
  wire  RVCExpander_1_io_rvc;
  wire [1:0] T_497;
  wire  T_498;
  wire  T_500;
  wire [3:0] T_501;
  wire  T_502;
  wire [1:0] T_504;
  wire  T_505;
  wire [1:0] T_506;
  wire  T_507;
  wire  T_508;
  wire  T_509;
  wire  T_510;
  wire [1:0] T_511;
  wire  T_512;
  wire [1:0] T_516;
  wire  T_517;
  wire  T_518;
  wire [1:0] T_522;
  wire  T_523;
  wire  T_524;
  wire  T_525;
  wire  T_526;
  wire [1:0] T_527;
  wire  T_528;
  wire  T_536;
  wire [3:0] T_544;
  wire  T_545;
  wire  T_546;
  wire  T_547;
  wire  T_548;
  wire [2:0] T_553;
  wire [1:0] T_554;
  wire [1:0] T_555;
  wire [1:0] GEN_30;
  RVCExpander RVCExpander_1 (
    .clk(RVCExpander_1_clk),
    .reset(RVCExpander_1_reset),
    .io_in(RVCExpander_1_io_in),
    .io_out_bits(RVCExpander_1_io_out_bits),
    .io_out_rd(RVCExpander_1_io_out_rd),
    .io_out_rs1(RVCExpander_1_io_out_rs1),
    .io_out_rs2(RVCExpander_1_io_out_rs2),
    .io_out_rs3(RVCExpander_1_io_out_rs3),
    .io_rvc(RVCExpander_1_io_rvc)
  );
  assign io_imem_ready = T_392;
  assign io_pc = T_495;
  assign io_btb_resp_taken = T_484_taken;
  assign io_btb_resp_mask = T_484_mask;
  assign io_btb_resp_bridx = T_484_bridx;
  assign io_btb_resp_target = T_484_target;
  assign io_btb_resp_entry = T_484_entry;
  assign io_btb_resp_bht_history = T_484_bht_history;
  assign io_btb_resp_bht_value = T_484_bht_value;
  assign io_inst_0_valid = T_526;
  assign io_inst_0_bits_pf0 = T_528;
  assign io_inst_0_bits_pf1 = T_536;
  assign io_inst_0_bits_replay = T_510;
  assign io_inst_0_bits_btb_hit = T_547;
  assign io_inst_0_bits_rvc = RVCExpander_1_io_rvc;
  assign io_inst_0_bits_inst_bits = RVCExpander_1_io_out_bits;
  assign io_inst_0_bits_inst_rd = RVCExpander_1_io_out_rd;
  assign io_inst_0_bits_inst_rs1 = RVCExpander_1_io_out_rs1;
  assign io_inst_0_bits_inst_rs2 = RVCExpander_1_io_out_rs2;
  assign io_inst_0_bits_inst_rs3 = RVCExpander_1_io_out_rs3;
  assign pcWordBits = io_imem_bits_pc[1];
  assign nReady = GEN_30;
  assign T_375 = io_imem_bits_btb_valid & io_imem_bits_btb_bits_taken;
  assign T_377 = io_imem_bits_btb_bits_bridx + 1'h1;
  assign T_379 = T_375 ? T_377 : 2'h2;
  assign GEN_31 = {{1'd0}, pcWordBits};
  assign T_380 = T_379 - GEN_31;
  assign nIC = T_380[1:0];
  assign GEN_32 = {{1'd0}, nBufValid};
  assign T_381 = nReady - GEN_32;
  assign nICReady = T_381[1:0];
  assign T_383 = io_imem_valid ? nIC : 2'h0;
  assign T_384 = T_383 + GEN_32;
  assign nValid = T_384[1:0];
  assign T_385 = nReady >= GEN_32;
  assign T_386 = nICReady >= nIC;
  assign T_388 = nIC - nICReady;
  assign T_389 = T_388[1:0];
  assign T_390 = 2'h1 >= T_389;
  assign T_391 = T_386 | T_390;
  assign T_392 = T_385 & T_391;
  assign T_395 = GEN_32 - nReady;
  assign T_396 = T_395[1:0];
  assign T_397 = T_385 ? 2'h0 : T_396;
  assign T_399 = io_imem_valid & T_385;
  assign T_400 = nICReady < nIC;
  assign T_401 = T_399 & T_400;
  assign T_406 = T_401 & T_390;
  assign T_407 = GEN_31 + nICReady;
  assign T_408 = T_407[1:0];
  assign T_411 = io_imem_bits_data[31:16];
  assign T_412 = {T_411,T_411};
  assign T_413 = {T_412,io_imem_bits_data};
  assign GEN_39 = {{4'd0}, T_408};
  assign T_414 = GEN_39 << 4;
  assign T_415 = T_413 >> T_414;
  assign T_416 = T_415[15:0];
  assign T_418 = io_imem_bits_pc & 40'hfffffffffc;
  assign GEN_40 = {{1'd0}, nICReady};
  assign T_419 = GEN_40 << 1;
  assign GEN_41 = {{37'd0}, T_419};
  assign T_420 = io_imem_bits_pc + GEN_41;
  assign T_421 = T_420[39:0];
  assign T_422 = T_421 & 40'h3;
  assign T_423 = T_418 | T_422;
  assign GEN_42 = {{1'd0}, io_imem_bits_btb_bits_bridx};
  assign T_424 = GEN_42 + nICReady;
  assign T_425 = T_424[1:0];
  assign GEN_0 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_taken : ibufBTBResp_taken;
  assign GEN_1 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_mask : ibufBTBResp_mask;
  assign GEN_2 = io_imem_bits_btb_valid ? T_425 : {{1'd0}, ibufBTBResp_bridx};
  assign GEN_3 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_target : ibufBTBResp_target;
  assign GEN_4 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_entry : ibufBTBResp_entry;
  assign GEN_5 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_bht_history : ibufBTBResp_bht_history;
  assign GEN_6 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_bht_value : ibufBTBResp_bht_value;
  assign GEN_7 = T_406 ? T_389 : T_397;
  assign GEN_8 = T_406 ? io_imem_bits_btb_valid : buf_btb_valid;
  assign GEN_9 = T_406 ? io_imem_bits_btb_bits_taken : buf_btb_bits_taken;
  assign GEN_10 = T_406 ? io_imem_bits_btb_bits_mask : buf_btb_bits_mask;
  assign GEN_11 = T_406 ? io_imem_bits_btb_bits_bridx : buf_btb_bits_bridx;
  assign GEN_12 = T_406 ? io_imem_bits_btb_bits_target : buf_btb_bits_target;
  assign GEN_13 = T_406 ? io_imem_bits_btb_bits_entry : buf_btb_bits_entry;
  assign GEN_14 = T_406 ? io_imem_bits_btb_bits_bht_history : buf_btb_bits_bht_history;
  assign GEN_15 = T_406 ? io_imem_bits_btb_bits_bht_value : buf_btb_bits_bht_value;
  assign GEN_16 = T_406 ? T_423 : buf_pc;
  assign GEN_17 = T_406 ? {{16'd0}, T_416} : buf_data;
  assign GEN_18 = T_406 ? io_imem_bits_mask : buf_mask;
  assign GEN_19 = T_406 ? io_imem_bits_xcpt_if : buf_xcpt_if;
  assign GEN_20 = T_406 ? io_imem_bits_replay : buf_replay;
  assign GEN_21 = T_406 ? io_imem_bits_btb_valid : ibufBTBHit;
  assign GEN_22 = T_406 ? GEN_0 : ibufBTBResp_taken;
  assign GEN_23 = T_406 ? GEN_1 : ibufBTBResp_mask;
  assign GEN_24 = T_406 ? GEN_2 : {{1'd0}, ibufBTBResp_bridx};
  assign GEN_25 = T_406 ? GEN_3 : ibufBTBResp_target;
  assign GEN_26 = T_406 ? GEN_4 : ibufBTBResp_entry;
  assign GEN_27 = T_406 ? GEN_5 : ibufBTBResp_bht_history;
  assign GEN_28 = T_406 ? GEN_6 : ibufBTBResp_bht_value;
  assign GEN_29 = io_kill ? 2'h0 : GEN_7;
  assign T_428 = 2'h2 + GEN_32;
  assign T_429 = T_428[1:0];
  assign T_430 = T_429 - GEN_31;
  assign T_431 = T_430[1:0];
  assign T_432 = io_imem_bits_data[15:0];
  assign T_433 = {T_432,T_432};
  assign T_434 = {io_imem_bits_data,T_433};
  assign T_435 = T_434[63:48];
  assign T_436 = {T_435,T_435};
  assign T_437 = {T_436,T_436};
  assign T_438 = {T_437,T_434};
  assign GEN_45 = {{4'd0}, T_431};
  assign T_439 = GEN_45 << 4;
  assign GEN_46 = {{63'd0}, T_438};
  assign T_440 = GEN_46 << T_439;
  assign icData = T_440[95:64];
  assign GEN_47 = {{4'd0}, nBufValid};
  assign T_443 = GEN_47 << 4;
  assign T_444 = 63'hffffffff << T_443;
  assign icMask = T_444[31:0];
  assign T_445 = icData & icMask;
  assign T_446 = ~ icMask;
  assign T_447 = buf_data & T_446;
  assign inst = T_445 | T_447;
  assign T_449 = 4'h1 << nValid;
  assign T_451 = T_449 - 4'h1;
  assign T_452 = T_451[3:0];
  assign valid = T_452[1:0];
  assign T_454 = 2'h1 << nBufValid;
  assign T_456 = T_454 - 2'h1;
  assign bufMask = T_456[1:0];
  assign T_458 = buf_xcpt_if ? bufMask : 2'h0;
  assign T_459 = ~ bufMask;
  assign T_461 = io_imem_bits_xcpt_if ? T_459 : 2'h0;
  assign T_462 = T_458 | T_461;
  assign xcpt_if = valid & T_462;
  assign T_464 = buf_replay ? bufMask : 2'h0;
  assign T_467 = io_imem_bits_replay ? T_459 : 2'h0;
  assign T_468 = T_464 | T_467;
  assign ic_replay = valid & T_468;
  assign T_470 = 2'h1 << ibufBTBResp_bridx;
  assign ibufBTBHitMask = ibufBTBHit ? T_470 : 2'h0;
  assign T_472 = io_imem_bits_btb_bits_bridx + nBufValid;
  assign T_473 = T_472 - GEN_31;
  assign T_474 = T_473[1:0];
  assign T_476 = 4'h1 << T_474;
  assign icBTBHitMask = io_imem_bits_btb_valid ? T_476 : 4'h0;
  assign T_478 = ibufBTBHitMask & bufMask;
  assign GEN_49 = {{2'd0}, T_459};
  assign T_480 = icBTBHitMask & GEN_49;
  assign GEN_50 = {{2'd0}, T_478};
  assign btbHitMask = GEN_50 | T_480;
  assign T_483 = T_478 != 2'h0;
  assign T_484_taken = T_483 ? ibufBTBResp_taken : io_imem_bits_btb_bits_taken;
  assign T_484_mask = T_483 ? ibufBTBResp_mask : io_imem_bits_btb_bits_mask;
  assign T_484_bridx = T_483 ? ibufBTBResp_bridx : io_imem_bits_btb_bits_bridx;
  assign T_484_target = T_483 ? ibufBTBResp_target : io_imem_bits_btb_bits_target;
  assign T_484_entry = T_483 ? ibufBTBResp_entry : io_imem_bits_btb_bits_entry;
  assign T_484_bht_history = T_483 ? ibufBTBResp_bht_history : io_imem_bits_btb_bits_bht_history;
  assign T_484_bht_value = T_483 ? ibufBTBResp_bht_value : io_imem_bits_btb_bits_bht_value;
  assign T_494 = nBufValid > 1'h0;
  assign T_495 = T_494 ? buf_pc : io_imem_bits_pc;
  assign RVCExpander_1_clk = clk;
  assign RVCExpander_1_reset = reset;
  assign RVCExpander_1_io_in = inst;
  assign T_497 = ic_replay >> 1'h0;
  assign T_498 = T_497[0];
  assign T_500 = RVCExpander_1_io_rvc == 1'h0;
  assign T_501 = btbHitMask >> 1'h0;
  assign T_502 = T_501[0];
  assign T_504 = 1'h0 + 1'h1;
  assign T_505 = T_504[0:0];
  assign T_506 = ic_replay >> T_505;
  assign T_507 = T_506[0];
  assign T_508 = T_502 | T_507;
  assign T_509 = T_500 & T_508;
  assign T_510 = T_498 | T_509;
  assign T_511 = valid >> 1'h0;
  assign T_512 = T_511[0];
  assign T_516 = valid >> T_505;
  assign T_517 = T_516[0];
  assign T_518 = RVCExpander_1_io_rvc | T_517;
  assign T_522 = xcpt_if >> T_505;
  assign T_523 = T_522[0];
  assign T_524 = T_518 | T_523;
  assign T_525 = T_524 | T_510;
  assign T_526 = T_512 & T_525;
  assign T_527 = xcpt_if >> 1'h0;
  assign T_528 = T_527[0];
  assign T_536 = T_500 & T_523;
  assign T_544 = btbHitMask >> T_505;
  assign T_545 = T_544[0];
  assign T_546 = T_500 & T_545;
  assign T_547 = T_502 | T_546;
  assign T_548 = io_inst_0_ready & io_inst_0_valid;
  assign T_553 = 2'h0 + 2'h2;
  assign T_554 = T_553[1:0];
  assign T_555 = RVCExpander_1_io_rvc ? {{1'd0}, T_505} : T_554;
  assign GEN_30 = T_548 ? T_555 : 2'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  nBufValid = GEN_33[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  buf_btb_valid = GEN_34[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {1{$random}};
  buf_btb_bits_taken = GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  buf_btb_bits_mask = GEN_36[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  buf_btb_bits_bridx = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {2{$random}};
  buf_btb_bits_target = GEN_38[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  buf_btb_bits_entry = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  buf_btb_bits_bht_history = GEN_44[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  buf_btb_bits_bht_value = GEN_48[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {2{$random}};
  buf_pc = GEN_51[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  buf_data = GEN_52[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {1{$random}};
  buf_mask = GEN_53[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {1{$random}};
  buf_xcpt_if = GEN_54[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {1{$random}};
  buf_replay = GEN_55[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {1{$random}};
  ibufBTBHit = GEN_56[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {1{$random}};
  ibufBTBResp_taken = GEN_57[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_58 = {1{$random}};
  ibufBTBResp_mask = GEN_58[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_59 = {1{$random}};
  ibufBTBResp_bridx = GEN_59[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_60 = {2{$random}};
  ibufBTBResp_target = GEN_60[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_61 = {1{$random}};
  ibufBTBResp_entry = GEN_61[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_62 = {1{$random}};
  ibufBTBResp_bht_history = GEN_62[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_63 = {1{$random}};
  ibufBTBResp_bht_value = GEN_63[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      nBufValid <= 1'h0;
    end else begin
      nBufValid <= GEN_29[0];
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_valid <= io_imem_bits_btb_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_taken <= io_imem_bits_btb_bits_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_mask <= io_imem_bits_btb_bits_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_bridx <= io_imem_bits_btb_bits_bridx;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_target <= io_imem_bits_btb_bits_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_entry <= io_imem_bits_btb_bits_entry;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_bht_history <= io_imem_bits_btb_bits_bht_history;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_bht_value <= io_imem_bits_btb_bits_bht_value;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_pc <= T_423;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_data <= {{16'd0}, T_416};
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_mask <= io_imem_bits_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_xcpt_if <= io_imem_bits_xcpt_if;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_replay <= io_imem_bits_replay;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        ibufBTBHit <= io_imem_bits_btb_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_taken <= io_imem_bits_btb_bits_taken;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_mask <= io_imem_bits_btb_bits_mask;
        end
      end
    end
    if(1'h0) begin
    end else begin
      ibufBTBResp_bridx <= GEN_24[0];
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_target <= io_imem_bits_btb_bits_target;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_entry <= io_imem_bits_btb_bits_entry;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_bht_history <= io_imem_bits_btb_bits_bht_history;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_bht_value <= io_imem_bits_btb_bits_bht_value;
        end
      end
    end
  end
endmodule
module CSRFile(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip,
  input  [11:0] io_rw_addr,
  input  [2:0] io_rw_cmd,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  output  io_csr_stall,
  output  io_csr_xcpt,
  output  io_eret,
  output  io_singleStep,
  output  io_status_debug,
  output [1:0] io_status_prv,
  output  io_status_sd,
  output [30:0] io_status_zero3,
  output  io_status_sd_rv32,
  output [1:0] io_status_zero2,
  output [4:0] io_status_vm,
  output [3:0] io_status_zero1,
  output  io_status_mxr,
  output  io_status_pum,
  output  io_status_mprv,
  output [1:0] io_status_xs,
  output [1:0] io_status_fs,
  output [1:0] io_status_mpp,
  output [1:0] io_status_hpp,
  output  io_status_spp,
  output  io_status_mpie,
  output  io_status_hpie,
  output  io_status_spie,
  output  io_status_upie,
  output  io_status_mie,
  output  io_status_hie,
  output  io_status_sie,
  output  io_status_uie,
  output [6:0] io_ptbr_asid,
  output [37:0] io_ptbr_ppn,
  output [39:0] io_evec,
  input   io_exception,
  input   io_retire,
  input  [63:0] io_cause,
  input  [39:0] io_pc,
  input  [39:0] io_badaddr,
  output  io_fatc,
  output [63:0] io_time,
  output [2:0] io_fcsr_rm,
  input   io_fcsr_flags_valid,
  input  [4:0] io_fcsr_flags_bits,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [63:0] io_rocc_cmd_bits_rs1,
  output [63:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_cmd_bits_status_debug,
  output [1:0] io_rocc_cmd_bits_status_prv,
  output  io_rocc_cmd_bits_status_sd,
  output [30:0] io_rocc_cmd_bits_status_zero3,
  output  io_rocc_cmd_bits_status_sd_rv32,
  output [1:0] io_rocc_cmd_bits_status_zero2,
  output [4:0] io_rocc_cmd_bits_status_vm,
  output [3:0] io_rocc_cmd_bits_status_zero1,
  output  io_rocc_cmd_bits_status_mxr,
  output  io_rocc_cmd_bits_status_pum,
  output  io_rocc_cmd_bits_status_mprv,
  output [1:0] io_rocc_cmd_bits_status_xs,
  output [1:0] io_rocc_cmd_bits_status_fs,
  output [1:0] io_rocc_cmd_bits_status_mpp,
  output [1:0] io_rocc_cmd_bits_status_hpp,
  output  io_rocc_cmd_bits_status_spp,
  output  io_rocc_cmd_bits_status_mpie,
  output  io_rocc_cmd_bits_status_hpie,
  output  io_rocc_cmd_bits_status_spie,
  output  io_rocc_cmd_bits_status_upie,
  output  io_rocc_cmd_bits_status_mie,
  output  io_rocc_cmd_bits_status_hie,
  output  io_rocc_cmd_bits_status_sie,
  output  io_rocc_cmd_bits_status_uie,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [63:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [39:0] io_rocc_mem_req_bits_addr,
  input  [5:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [63:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [63:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [39:0] io_rocc_mem_resp_bits_addr,
  output [5:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [63:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [63:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [63:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input   io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [10:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output  io_rocc_autl_grant_bits_client_xact_id,
  output [1:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception,
  output  io_interrupt,
  output [63:0] io_interrupt_cause,
  output [3:0] io_bp_0_control_ttype,
  output  io_bp_0_control_dmode,
  output [5:0] io_bp_0_control_maskmax,
  output [39:0] io_bp_0_control_reserved,
  output  io_bp_0_control_action,
  output  io_bp_0_control_chain,
  output [1:0] io_bp_0_control_zero,
  output [1:0] io_bp_0_control_tmatch,
  output  io_bp_0_control_m,
  output  io_bp_0_control_h,
  output  io_bp_0_control_s,
  output  io_bp_0_control_u,
  output  io_bp_0_control_x,
  output  io_bp_0_control_w,
  output  io_bp_0_control_r,
  output [38:0] io_bp_0_address
);
  wire  T_4982_debug;
  wire [1:0] T_4982_prv;
  wire  T_4982_sd;
  wire [30:0] T_4982_zero3;
  wire  T_4982_sd_rv32;
  wire [1:0] T_4982_zero2;
  wire [4:0] T_4982_vm;
  wire [3:0] T_4982_zero1;
  wire  T_4982_mxr;
  wire  T_4982_pum;
  wire  T_4982_mprv;
  wire [1:0] T_4982_xs;
  wire [1:0] T_4982_fs;
  wire [1:0] T_4982_mpp;
  wire [1:0] T_4982_hpp;
  wire  T_4982_spp;
  wire  T_4982_mpie;
  wire  T_4982_hpie;
  wire  T_4982_spie;
  wire  T_4982_upie;
  wire  T_4982_mie;
  wire  T_4982_hie;
  wire  T_4982_sie;
  wire  T_4982_uie;
  wire [66:0] T_5008;
  wire  T_5009;
  wire  T_5010;
  wire  T_5011;
  wire  T_5012;
  wire  T_5013;
  wire  T_5014;
  wire  T_5015;
  wire  T_5016;
  wire  T_5017;
  wire [1:0] T_5018;
  wire [1:0] T_5019;
  wire [1:0] T_5020;
  wire [1:0] T_5021;
  wire  T_5022;
  wire  T_5023;
  wire  T_5024;
  wire [3:0] T_5025;
  wire [4:0] T_5026;
  wire [1:0] T_5027;
  wire  T_5028;
  wire [30:0] T_5029;
  wire  T_5030;
  wire [1:0] T_5031;
  wire  T_5032;
  wire  reset_mstatus_debug;
  wire [1:0] reset_mstatus_prv;
  wire  reset_mstatus_sd;
  wire [30:0] reset_mstatus_zero3;
  wire  reset_mstatus_sd_rv32;
  wire [1:0] reset_mstatus_zero2;
  wire [4:0] reset_mstatus_vm;
  wire [3:0] reset_mstatus_zero1;
  wire  reset_mstatus_mxr;
  wire  reset_mstatus_pum;
  wire  reset_mstatus_mprv;
  wire [1:0] reset_mstatus_xs;
  wire [1:0] reset_mstatus_fs;
  wire [1:0] reset_mstatus_mpp;
  wire [1:0] reset_mstatus_hpp;
  wire  reset_mstatus_spp;
  wire  reset_mstatus_mpie;
  wire  reset_mstatus_hpie;
  wire  reset_mstatus_spie;
  wire  reset_mstatus_upie;
  wire  reset_mstatus_mie;
  wire  reset_mstatus_hie;
  wire  reset_mstatus_sie;
  wire  reset_mstatus_uie;
  reg  reg_mstatus_debug;
  reg [31:0] GEN_120;
  reg [1:0] reg_mstatus_prv;
  reg [31:0] GEN_121;
  reg  reg_mstatus_sd;
  reg [31:0] GEN_122;
  reg [30:0] reg_mstatus_zero3;
  reg [31:0] GEN_123;
  reg  reg_mstatus_sd_rv32;
  reg [31:0] GEN_124;
  reg [1:0] reg_mstatus_zero2;
  reg [31:0] GEN_125;
  reg [4:0] reg_mstatus_vm;
  reg [31:0] GEN_126;
  reg [3:0] reg_mstatus_zero1;
  reg [31:0] GEN_127;
  reg  reg_mstatus_mxr;
  reg [31:0] GEN_128;
  reg  reg_mstatus_pum;
  reg [31:0] GEN_129;
  reg  reg_mstatus_mprv;
  reg [31:0] GEN_130;
  reg [1:0] reg_mstatus_xs;
  reg [31:0] GEN_131;
  reg [1:0] reg_mstatus_fs;
  reg [31:0] GEN_132;
  reg [1:0] reg_mstatus_mpp;
  reg [31:0] GEN_133;
  reg [1:0] reg_mstatus_hpp;
  reg [31:0] GEN_134;
  reg  reg_mstatus_spp;
  reg [31:0] GEN_135;
  reg  reg_mstatus_mpie;
  reg [31:0] GEN_136;
  reg  reg_mstatus_hpie;
  reg [31:0] GEN_137;
  reg  reg_mstatus_spie;
  reg [31:0] GEN_138;
  reg  reg_mstatus_upie;
  reg [31:0] GEN_139;
  reg  reg_mstatus_mie;
  reg [31:0] GEN_140;
  reg  reg_mstatus_hie;
  reg [31:0] GEN_141;
  reg  reg_mstatus_sie;
  reg [31:0] GEN_142;
  reg  reg_mstatus_uie;
  reg [31:0] GEN_143;
  wire [1:0] new_prv;
  wire [1:0] T_5121_xdebugver;
  wire  T_5121_ndreset;
  wire  T_5121_fullreset;
  wire [11:0] T_5121_zero3;
  wire  T_5121_ebreakm;
  wire  T_5121_ebreakh;
  wire  T_5121_ebreaks;
  wire  T_5121_ebreaku;
  wire  T_5121_zero2;
  wire  T_5121_stopcycle;
  wire  T_5121_stoptime;
  wire [2:0] T_5121_cause;
  wire  T_5121_debugint;
  wire  T_5121_zero1;
  wire  T_5121_halt;
  wire  T_5121_step;
  wire [1:0] T_5121_prv;
  wire [31:0] T_5140;
  wire [1:0] T_5141;
  wire  T_5142;
  wire  T_5143;
  wire  T_5144;
  wire  T_5145;
  wire [2:0] T_5146;
  wire  T_5147;
  wire  T_5148;
  wire  T_5149;
  wire  T_5150;
  wire  T_5151;
  wire  T_5152;
  wire  T_5153;
  wire [11:0] T_5154;
  wire  T_5155;
  wire  T_5156;
  wire [1:0] T_5157;
  wire [1:0] reset_dcsr_xdebugver;
  wire  reset_dcsr_ndreset;
  wire  reset_dcsr_fullreset;
  wire [11:0] reset_dcsr_zero3;
  wire  reset_dcsr_ebreakm;
  wire  reset_dcsr_ebreakh;
  wire  reset_dcsr_ebreaks;
  wire  reset_dcsr_ebreaku;
  wire  reset_dcsr_zero2;
  wire  reset_dcsr_stopcycle;
  wire  reset_dcsr_stoptime;
  wire [2:0] reset_dcsr_cause;
  wire  reset_dcsr_debugint;
  wire  reset_dcsr_zero1;
  wire  reset_dcsr_halt;
  wire  reset_dcsr_step;
  wire [1:0] reset_dcsr_prv;
  reg [1:0] reg_dcsr_xdebugver;
  reg [31:0] GEN_144;
  reg  reg_dcsr_ndreset;
  reg [31:0] GEN_145;
  reg  reg_dcsr_fullreset;
  reg [31:0] GEN_146;
  reg [11:0] reg_dcsr_zero3;
  reg [31:0] GEN_147;
  reg  reg_dcsr_ebreakm;
  reg [31:0] GEN_148;
  reg  reg_dcsr_ebreakh;
  reg [31:0] GEN_149;
  reg  reg_dcsr_ebreaks;
  reg [31:0] GEN_150;
  reg  reg_dcsr_ebreaku;
  reg [31:0] GEN_151;
  reg  reg_dcsr_zero2;
  reg [31:0] GEN_152;
  reg  reg_dcsr_stopcycle;
  reg [31:0] GEN_153;
  reg  reg_dcsr_stoptime;
  reg [31:0] GEN_154;
  reg [2:0] reg_dcsr_cause;
  reg [31:0] GEN_155;
  reg  reg_dcsr_debugint;
  reg [31:0] GEN_156;
  reg  reg_dcsr_zero1;
  reg [31:0] GEN_157;
  reg  reg_dcsr_halt;
  reg [31:0] GEN_158;
  reg  reg_dcsr_step;
  reg [31:0] GEN_159;
  reg [1:0] reg_dcsr_prv;
  reg [31:0] GEN_160;
  wire  T_5223_rocc;
  wire  T_5223_meip;
  wire  T_5223_heip;
  wire  T_5223_seip;
  wire  T_5223_ueip;
  wire  T_5223_mtip;
  wire  T_5223_htip;
  wire  T_5223_stip;
  wire  T_5223_utip;
  wire  T_5223_msip;
  wire  T_5223_hsip;
  wire  T_5223_ssip;
  wire  T_5223_usip;
  wire [12:0] T_5238;
  wire  T_5239;
  wire  T_5240;
  wire  T_5241;
  wire  T_5242;
  wire  T_5243;
  wire  T_5244;
  wire  T_5245;
  wire  T_5246;
  wire  T_5247;
  wire  T_5248;
  wire  T_5249;
  wire  T_5250;
  wire  T_5251;
  wire  T_5252_rocc;
  wire  T_5252_meip;
  wire  T_5252_heip;
  wire  T_5252_seip;
  wire  T_5252_ueip;
  wire  T_5252_mtip;
  wire  T_5252_htip;
  wire  T_5252_stip;
  wire  T_5252_utip;
  wire  T_5252_msip;
  wire  T_5252_hsip;
  wire  T_5252_ssip;
  wire  T_5252_usip;
  wire  T_5273_rocc;
  wire  T_5273_meip;
  wire  T_5273_heip;
  wire  T_5273_seip;
  wire  T_5273_ueip;
  wire  T_5273_mtip;
  wire  T_5273_htip;
  wire  T_5273_stip;
  wire  T_5273_utip;
  wire  T_5273_msip;
  wire  T_5273_hsip;
  wire  T_5273_ssip;
  wire  T_5273_usip;
  wire [1:0] T_5290;
  wire [2:0] T_5291;
  wire [1:0] T_5292;
  wire [2:0] T_5293;
  wire [5:0] T_5294;
  wire [1:0] T_5295;
  wire [2:0] T_5296;
  wire [1:0] T_5297;
  wire [1:0] T_5298;
  wire [3:0] T_5299;
  wire [6:0] T_5300;
  wire [12:0] supported_interrupts;
  wire  exception;
  reg  reg_debug;
  reg [31:0] GEN_161;
  reg [39:0] reg_dpc;
  reg [63:0] GEN_162;
  reg [63:0] reg_dscratch;
  reg [63:0] GEN_163;
  reg  reg_singleStepped;
  reg [31:0] GEN_164;
  wire  T_5317;
  wire  GEN_36;
  wire  T_5320;
  wire  GEN_37;
  wire  T_5331;
  wire  T_5333;
  wire  T_5334;
  wire  T_5335;
  wire  T_5337;
  reg  reg_tselect;
  reg [31:0] GEN_165;
  reg [3:0] reg_bp_0_control_ttype;
  reg [31:0] GEN_166;
  reg  reg_bp_0_control_dmode;
  reg [31:0] GEN_167;
  reg [5:0] reg_bp_0_control_maskmax;
  reg [31:0] GEN_168;
  reg [39:0] reg_bp_0_control_reserved;
  reg [63:0] GEN_169;
  reg  reg_bp_0_control_action;
  reg [31:0] GEN_170;
  reg  reg_bp_0_control_chain;
  reg [31:0] GEN_171;
  reg [1:0] reg_bp_0_control_zero;
  reg [31:0] GEN_172;
  reg [1:0] reg_bp_0_control_tmatch;
  reg [31:0] GEN_173;
  reg  reg_bp_0_control_m;
  reg [31:0] GEN_174;
  reg  reg_bp_0_control_h;
  reg [31:0] GEN_175;
  reg  reg_bp_0_control_s;
  reg [31:0] GEN_176;
  reg  reg_bp_0_control_u;
  reg [31:0] GEN_177;
  reg  reg_bp_0_control_x;
  reg [31:0] GEN_178;
  reg  reg_bp_0_control_w;
  reg [31:0] GEN_179;
  reg  reg_bp_0_control_r;
  reg [31:0] GEN_180;
  reg [38:0] reg_bp_0_address;
  reg [63:0] GEN_181;
  reg [3:0] reg_bp_1_control_ttype;
  reg [31:0] GEN_182;
  reg  reg_bp_1_control_dmode;
  reg [31:0] GEN_183;
  reg [5:0] reg_bp_1_control_maskmax;
  reg [31:0] GEN_184;
  reg [39:0] reg_bp_1_control_reserved;
  reg [63:0] GEN_185;
  reg  reg_bp_1_control_action;
  reg [31:0] GEN_186;
  reg  reg_bp_1_control_chain;
  reg [31:0] GEN_187;
  reg [1:0] reg_bp_1_control_zero;
  reg [31:0] GEN_188;
  reg [1:0] reg_bp_1_control_tmatch;
  reg [31:0] GEN_189;
  reg  reg_bp_1_control_m;
  reg [31:0] GEN_190;
  reg  reg_bp_1_control_h;
  reg [31:0] GEN_191;
  reg  reg_bp_1_control_s;
  reg [31:0] GEN_192;
  reg  reg_bp_1_control_u;
  reg [31:0] GEN_193;
  reg  reg_bp_1_control_x;
  reg [31:0] GEN_194;
  reg  reg_bp_1_control_w;
  reg [31:0] GEN_195;
  reg  reg_bp_1_control_r;
  reg [31:0] GEN_196;
  reg [38:0] reg_bp_1_address;
  reg [63:0] GEN_197;
  reg [63:0] reg_mie;
  reg [63:0] GEN_198;
  reg [63:0] reg_mideleg;
  reg [63:0] GEN_199;
  reg [63:0] reg_medeleg;
  reg [63:0] GEN_200;
  reg  reg_mip_rocc;
  reg [31:0] GEN_201;
  reg  reg_mip_meip;
  reg [31:0] GEN_202;
  reg  reg_mip_heip;
  reg [31:0] GEN_203;
  reg  reg_mip_seip;
  reg [31:0] GEN_204;
  reg  reg_mip_ueip;
  reg [31:0] GEN_205;
  reg  reg_mip_mtip;
  reg [31:0] GEN_206;
  reg  reg_mip_htip;
  reg [31:0] GEN_207;
  reg  reg_mip_stip;
  reg [31:0] GEN_208;
  reg  reg_mip_utip;
  reg [31:0] GEN_209;
  reg  reg_mip_msip;
  reg [31:0] GEN_210;
  reg  reg_mip_hsip;
  reg [31:0] GEN_211;
  reg  reg_mip_ssip;
  reg [31:0] GEN_212;
  reg  reg_mip_usip;
  reg [31:0] GEN_213;
  reg [39:0] reg_mepc;
  reg [63:0] GEN_214;
  reg [63:0] reg_mcause;
  reg [63:0] GEN_215;
  reg [39:0] reg_mbadaddr;
  reg [63:0] GEN_216;
  reg [63:0] reg_mscratch;
  reg [63:0] GEN_217;
  reg [31:0] reg_mtvec;
  reg [31:0] GEN_218;
  reg [31:0] reg_mucounteren;
  reg [31:0] GEN_219;
  reg [31:0] reg_mscounteren;
  reg [31:0] GEN_220;
  reg [39:0] reg_sepc;
  reg [63:0] GEN_221;
  reg [63:0] reg_scause;
  reg [63:0] GEN_222;
  reg [39:0] reg_sbadaddr;
  reg [63:0] GEN_223;
  reg [63:0] reg_sscratch;
  reg [63:0] GEN_224;
  reg [38:0] reg_stvec;
  reg [63:0] GEN_225;
  reg [6:0] reg_sptbr_asid;
  reg [31:0] GEN_226;
  reg [37:0] reg_sptbr_ppn;
  reg [63:0] GEN_227;
  reg  reg_wfi;
  reg [31:0] GEN_228;
  reg [4:0] reg_fflags;
  reg [31:0] GEN_229;
  reg [2:0] reg_frm;
  reg [31:0] GEN_230;
  reg [5:0] T_5567;
  reg [31:0] GEN_231;
  wire [5:0] GEN_0;
  wire [6:0] T_5568;
  reg [57:0] T_5570;
  reg [63:0] GEN_232;
  wire  T_5571;
  wire [58:0] T_5573;
  wire [57:0] T_5574;
  wire [57:0] GEN_38;
  wire [63:0] T_5575;
  reg [5:0] T_5578;
  reg [31:0] GEN_233;
  wire [6:0] T_5579;
  reg [57:0] T_5581;
  reg [63:0] GEN_234;
  wire  T_5582;
  wire [58:0] T_5584;
  wire [57:0] T_5585;
  wire [57:0] GEN_39;
  wire [63:0] T_5586;
  wire  mip_rocc;
  wire  mip_meip;
  wire  mip_heip;
  wire  mip_seip;
  wire  mip_ueip;
  wire  mip_mtip;
  wire  mip_htip;
  wire  mip_stip;
  wire  mip_utip;
  wire  mip_msip;
  wire  mip_hsip;
  wire  mip_ssip;
  wire  mip_usip;
  wire [1:0] T_5600;
  wire [2:0] T_5601;
  wire [1:0] T_5602;
  wire [2:0] T_5603;
  wire [5:0] T_5604;
  wire [1:0] T_5605;
  wire [2:0] T_5606;
  wire [1:0] T_5607;
  wire [1:0] T_5608;
  wire [3:0] T_5609;
  wire [6:0] T_5610;
  wire [12:0] T_5611;
  wire [12:0] read_mip;
  wire [63:0] GEN_1;
  wire [63:0] pending_interrupts;
  wire  T_5613;
  wire  T_5615;
  wire  T_5617;
  wire  T_5618;
  wire  T_5619;
  wire  T_5620;
  wire [63:0] T_5621;
  wire [63:0] T_5622;
  wire [63:0] m_interrupts;
  wire  T_5627;
  wire  T_5629;
  wire  T_5630;
  wire  T_5631;
  wire  T_5632;
  wire [63:0] T_5633;
  wire [63:0] s_interrupts;
  wire [63:0] all_interrupts;
  wire  T_5636;
  wire  T_5637;
  wire  T_5638;
  wire  T_5639;
  wire  T_5640;
  wire  T_5641;
  wire  T_5642;
  wire  T_5643;
  wire  T_5644;
  wire  T_5645;
  wire  T_5646;
  wire  T_5647;
  wire  T_5648;
  wire  T_5649;
  wire  T_5650;
  wire  T_5651;
  wire  T_5652;
  wire  T_5653;
  wire  T_5654;
  wire  T_5655;
  wire  T_5656;
  wire  T_5657;
  wire  T_5658;
  wire  T_5659;
  wire  T_5660;
  wire  T_5661;
  wire  T_5662;
  wire  T_5663;
  wire  T_5664;
  wire  T_5665;
  wire  T_5666;
  wire  T_5667;
  wire  T_5668;
  wire  T_5669;
  wire  T_5670;
  wire  T_5671;
  wire  T_5672;
  wire  T_5673;
  wire  T_5674;
  wire  T_5675;
  wire  T_5676;
  wire  T_5677;
  wire  T_5678;
  wire  T_5679;
  wire  T_5680;
  wire  T_5681;
  wire  T_5682;
  wire  T_5683;
  wire  T_5684;
  wire  T_5685;
  wire  T_5686;
  wire  T_5687;
  wire  T_5688;
  wire  T_5689;
  wire  T_5690;
  wire  T_5691;
  wire  T_5692;
  wire  T_5693;
  wire  T_5694;
  wire  T_5695;
  wire  T_5696;
  wire  T_5697;
  wire  T_5698;
  wire [5:0] T_5764;
  wire [5:0] T_5765;
  wire [5:0] T_5766;
  wire [5:0] T_5767;
  wire [5:0] T_5768;
  wire [5:0] T_5769;
  wire [5:0] T_5770;
  wire [5:0] T_5771;
  wire [5:0] T_5772;
  wire [5:0] T_5773;
  wire [5:0] T_5774;
  wire [5:0] T_5775;
  wire [5:0] T_5776;
  wire [5:0] T_5777;
  wire [5:0] T_5778;
  wire [5:0] T_5779;
  wire [5:0] T_5780;
  wire [5:0] T_5781;
  wire [5:0] T_5782;
  wire [5:0] T_5783;
  wire [5:0] T_5784;
  wire [5:0] T_5785;
  wire [5:0] T_5786;
  wire [5:0] T_5787;
  wire [5:0] T_5788;
  wire [5:0] T_5789;
  wire [5:0] T_5790;
  wire [5:0] T_5791;
  wire [5:0] T_5792;
  wire [5:0] T_5793;
  wire [5:0] T_5794;
  wire [5:0] T_5795;
  wire [5:0] T_5796;
  wire [5:0] T_5797;
  wire [5:0] T_5798;
  wire [5:0] T_5799;
  wire [5:0] T_5800;
  wire [5:0] T_5801;
  wire [5:0] T_5802;
  wire [5:0] T_5803;
  wire [5:0] T_5804;
  wire [5:0] T_5805;
  wire [5:0] T_5806;
  wire [5:0] T_5807;
  wire [5:0] T_5808;
  wire [5:0] T_5809;
  wire [5:0] T_5810;
  wire [5:0] T_5811;
  wire [5:0] T_5812;
  wire [5:0] T_5813;
  wire [5:0] T_5814;
  wire [5:0] T_5815;
  wire [5:0] T_5816;
  wire [5:0] T_5817;
  wire [5:0] T_5818;
  wire [5:0] T_5819;
  wire [5:0] T_5820;
  wire [5:0] T_5821;
  wire [5:0] T_5822;
  wire [5:0] T_5823;
  wire [5:0] T_5824;
  wire [5:0] T_5825;
  wire [5:0] T_5826;
  wire [63:0] GEN_2;
  wire [64:0] T_5827;
  wire [63:0] interruptCause;
  wire  T_5829;
  wire  T_5832;
  wire  T_5833;
  wire  T_5838;
  wire  GEN_40;
  wire [63:0] GEN_41;
  wire  system_insn;
  wire  T_5841;
  wire  T_5843;
  wire  cpu_ren;
  wire  T_5844;
  wire  cpu_wen;
  wire [1:0] T_5845;
  wire [2:0] T_5846;
  wire [1:0] T_5847;
  wire [2:0] T_5848;
  wire [5:0] T_5849;
  wire [1:0] T_5850;
  wire [2:0] T_5851;
  wire [3:0] T_5852;
  wire [5:0] T_5853;
  wire [8:0] T_5854;
  wire [14:0] T_5855;
  wire [1:0] T_5856;
  wire [3:0] T_5857;
  wire [8:0] T_5858;
  wire [9:0] T_5859;
  wire [13:0] T_5860;
  wire [31:0] T_5861;
  wire [33:0] T_5862;
  wire [2:0] T_5863;
  wire [3:0] T_5864;
  wire [37:0] T_5865;
  wire [51:0] T_5866;
  wire [66:0] T_5867;
  wire [63:0] read_mstatus;
  wire [3:0] GEN_0_control_ttype;
  wire  GEN_0_control_dmode;
  wire [5:0] GEN_0_control_maskmax;
  wire [39:0] GEN_0_control_reserved;
  wire  GEN_0_control_action;
  wire  GEN_0_control_chain;
  wire [1:0] GEN_0_control_zero;
  wire [1:0] GEN_0_control_tmatch;
  wire  GEN_0_control_m;
  wire  GEN_0_control_h;
  wire  GEN_0_control_s;
  wire  GEN_0_control_u;
  wire  GEN_0_control_x;
  wire  GEN_0_control_w;
  wire  GEN_0_control_r;
  wire [38:0] GEN_0_address;
  wire [3:0] GEN_42;
  wire  GEN_43;
  wire [5:0] GEN_44;
  wire [39:0] GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire [1:0] GEN_48;
  wire [1:0] GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire [38:0] GEN_57;
  wire [3:0] GEN_1_control_ttype;
  wire  GEN_1_control_dmode;
  wire [5:0] GEN_1_control_maskmax;
  wire [39:0] GEN_1_control_reserved;
  wire  GEN_1_control_action;
  wire  GEN_1_control_chain;
  wire [1:0] GEN_1_control_zero;
  wire [1:0] GEN_1_control_tmatch;
  wire  GEN_1_control_m;
  wire  GEN_1_control_h;
  wire  GEN_1_control_s;
  wire  GEN_1_control_u;
  wire  GEN_1_control_x;
  wire  GEN_1_control_w;
  wire  GEN_1_control_r;
  wire [38:0] GEN_1_address;
  wire [1:0] T_5885;
  wire [3:0] GEN_2_control_ttype;
  wire  GEN_2_control_dmode;
  wire [5:0] GEN_2_control_maskmax;
  wire [39:0] GEN_2_control_reserved;
  wire  GEN_2_control_action;
  wire  GEN_2_control_chain;
  wire [1:0] GEN_2_control_zero;
  wire [1:0] GEN_2_control_tmatch;
  wire  GEN_2_control_m;
  wire  GEN_2_control_h;
  wire  GEN_2_control_s;
  wire  GEN_2_control_u;
  wire  GEN_2_control_x;
  wire  GEN_2_control_w;
  wire  GEN_2_control_r;
  wire [38:0] GEN_2_address;
  wire [2:0] T_5886;
  wire [3:0] GEN_3_control_ttype;
  wire  GEN_3_control_dmode;
  wire [5:0] GEN_3_control_maskmax;
  wire [39:0] GEN_3_control_reserved;
  wire  GEN_3_control_action;
  wire  GEN_3_control_chain;
  wire [1:0] GEN_3_control_zero;
  wire [1:0] GEN_3_control_tmatch;
  wire  GEN_3_control_m;
  wire  GEN_3_control_h;
  wire  GEN_3_control_s;
  wire  GEN_3_control_u;
  wire  GEN_3_control_x;
  wire  GEN_3_control_w;
  wire  GEN_3_control_r;
  wire [38:0] GEN_3_address;
  wire [3:0] GEN_4_control_ttype;
  wire  GEN_4_control_dmode;
  wire [5:0] GEN_4_control_maskmax;
  wire [39:0] GEN_4_control_reserved;
  wire  GEN_4_control_action;
  wire  GEN_4_control_chain;
  wire [1:0] GEN_4_control_zero;
  wire [1:0] GEN_4_control_tmatch;
  wire  GEN_4_control_m;
  wire  GEN_4_control_h;
  wire  GEN_4_control_s;
  wire  GEN_4_control_u;
  wire  GEN_4_control_x;
  wire  GEN_4_control_w;
  wire  GEN_4_control_r;
  wire [38:0] GEN_4_address;
  wire [1:0] T_5887;
  wire [3:0] GEN_5_control_ttype;
  wire  GEN_5_control_dmode;
  wire [5:0] GEN_5_control_maskmax;
  wire [39:0] GEN_5_control_reserved;
  wire  GEN_5_control_action;
  wire  GEN_5_control_chain;
  wire [1:0] GEN_5_control_zero;
  wire [1:0] GEN_5_control_tmatch;
  wire  GEN_5_control_m;
  wire  GEN_5_control_h;
  wire  GEN_5_control_s;
  wire  GEN_5_control_u;
  wire  GEN_5_control_x;
  wire  GEN_5_control_w;
  wire  GEN_5_control_r;
  wire [38:0] GEN_5_address;
  wire [3:0] GEN_6_control_ttype;
  wire  GEN_6_control_dmode;
  wire [5:0] GEN_6_control_maskmax;
  wire [39:0] GEN_6_control_reserved;
  wire  GEN_6_control_action;
  wire  GEN_6_control_chain;
  wire [1:0] GEN_6_control_zero;
  wire [1:0] GEN_6_control_tmatch;
  wire  GEN_6_control_m;
  wire  GEN_6_control_h;
  wire  GEN_6_control_s;
  wire  GEN_6_control_u;
  wire  GEN_6_control_x;
  wire  GEN_6_control_w;
  wire  GEN_6_control_r;
  wire [38:0] GEN_6_address;
  wire [1:0] T_5888;
  wire [3:0] T_5889;
  wire [6:0] T_5890;
  wire [3:0] GEN_7_control_ttype;
  wire  GEN_7_control_dmode;
  wire [5:0] GEN_7_control_maskmax;
  wire [39:0] GEN_7_control_reserved;
  wire  GEN_7_control_action;
  wire  GEN_7_control_chain;
  wire [1:0] GEN_7_control_zero;
  wire [1:0] GEN_7_control_tmatch;
  wire  GEN_7_control_m;
  wire  GEN_7_control_h;
  wire  GEN_7_control_s;
  wire  GEN_7_control_u;
  wire  GEN_7_control_x;
  wire  GEN_7_control_w;
  wire  GEN_7_control_r;
  wire [38:0] GEN_7_address;
  wire [3:0] GEN_8_control_ttype;
  wire  GEN_8_control_dmode;
  wire [5:0] GEN_8_control_maskmax;
  wire [39:0] GEN_8_control_reserved;
  wire  GEN_8_control_action;
  wire  GEN_8_control_chain;
  wire [1:0] GEN_8_control_zero;
  wire [1:0] GEN_8_control_tmatch;
  wire  GEN_8_control_m;
  wire  GEN_8_control_h;
  wire  GEN_8_control_s;
  wire  GEN_8_control_u;
  wire  GEN_8_control_x;
  wire  GEN_8_control_w;
  wire  GEN_8_control_r;
  wire [38:0] GEN_8_address;
  wire [3:0] T_5891;
  wire [3:0] GEN_9_control_ttype;
  wire  GEN_9_control_dmode;
  wire [5:0] GEN_9_control_maskmax;
  wire [39:0] GEN_9_control_reserved;
  wire  GEN_9_control_action;
  wire  GEN_9_control_chain;
  wire [1:0] GEN_9_control_zero;
  wire [1:0] GEN_9_control_tmatch;
  wire  GEN_9_control_m;
  wire  GEN_9_control_h;
  wire  GEN_9_control_s;
  wire  GEN_9_control_u;
  wire  GEN_9_control_x;
  wire  GEN_9_control_w;
  wire  GEN_9_control_r;
  wire [38:0] GEN_9_address;
  wire [3:0] GEN_10_control_ttype;
  wire  GEN_10_control_dmode;
  wire [5:0] GEN_10_control_maskmax;
  wire [39:0] GEN_10_control_reserved;
  wire  GEN_10_control_action;
  wire  GEN_10_control_chain;
  wire [1:0] GEN_10_control_zero;
  wire [1:0] GEN_10_control_tmatch;
  wire  GEN_10_control_m;
  wire  GEN_10_control_h;
  wire  GEN_10_control_s;
  wire  GEN_10_control_u;
  wire  GEN_10_control_x;
  wire  GEN_10_control_w;
  wire  GEN_10_control_r;
  wire [38:0] GEN_10_address;
  wire [1:0] T_5892;
  wire [5:0] T_5893;
  wire [3:0] GEN_11_control_ttype;
  wire  GEN_11_control_dmode;
  wire [5:0] GEN_11_control_maskmax;
  wire [39:0] GEN_11_control_reserved;
  wire  GEN_11_control_action;
  wire  GEN_11_control_chain;
  wire [1:0] GEN_11_control_zero;
  wire [1:0] GEN_11_control_tmatch;
  wire  GEN_11_control_m;
  wire  GEN_11_control_h;
  wire  GEN_11_control_s;
  wire  GEN_11_control_u;
  wire  GEN_11_control_x;
  wire  GEN_11_control_w;
  wire  GEN_11_control_r;
  wire [38:0] GEN_11_address;
  wire [3:0] GEN_12_control_ttype;
  wire  GEN_12_control_dmode;
  wire [5:0] GEN_12_control_maskmax;
  wire [39:0] GEN_12_control_reserved;
  wire  GEN_12_control_action;
  wire  GEN_12_control_chain;
  wire [1:0] GEN_12_control_zero;
  wire [1:0] GEN_12_control_tmatch;
  wire  GEN_12_control_m;
  wire  GEN_12_control_h;
  wire  GEN_12_control_s;
  wire  GEN_12_control_u;
  wire  GEN_12_control_x;
  wire  GEN_12_control_w;
  wire  GEN_12_control_r;
  wire [38:0] GEN_12_address;
  wire [45:0] T_5894;
  wire [3:0] GEN_13_control_ttype;
  wire  GEN_13_control_dmode;
  wire [5:0] GEN_13_control_maskmax;
  wire [39:0] GEN_13_control_reserved;
  wire  GEN_13_control_action;
  wire  GEN_13_control_chain;
  wire [1:0] GEN_13_control_zero;
  wire [1:0] GEN_13_control_tmatch;
  wire  GEN_13_control_m;
  wire  GEN_13_control_h;
  wire  GEN_13_control_s;
  wire  GEN_13_control_u;
  wire  GEN_13_control_x;
  wire  GEN_13_control_w;
  wire  GEN_13_control_r;
  wire [38:0] GEN_13_address;
  wire [3:0] GEN_14_control_ttype;
  wire  GEN_14_control_dmode;
  wire [5:0] GEN_14_control_maskmax;
  wire [39:0] GEN_14_control_reserved;
  wire  GEN_14_control_action;
  wire  GEN_14_control_chain;
  wire [1:0] GEN_14_control_zero;
  wire [1:0] GEN_14_control_tmatch;
  wire  GEN_14_control_m;
  wire  GEN_14_control_h;
  wire  GEN_14_control_s;
  wire  GEN_14_control_u;
  wire  GEN_14_control_x;
  wire  GEN_14_control_w;
  wire  GEN_14_control_r;
  wire [38:0] GEN_14_address;
  wire [4:0] T_5895;
  wire [50:0] T_5896;
  wire [56:0] T_5897;
  wire [63:0] T_5898;
  wire [3:0] GEN_15_control_ttype;
  wire  GEN_15_control_dmode;
  wire [5:0] GEN_15_control_maskmax;
  wire [39:0] GEN_15_control_reserved;
  wire  GEN_15_control_action;
  wire  GEN_15_control_chain;
  wire [1:0] GEN_15_control_zero;
  wire [1:0] GEN_15_control_tmatch;
  wire  GEN_15_control_m;
  wire  GEN_15_control_h;
  wire  GEN_15_control_s;
  wire  GEN_15_control_u;
  wire  GEN_15_control_x;
  wire  GEN_15_control_w;
  wire  GEN_15_control_r;
  wire [38:0] GEN_15_address;
  wire  T_5916;
  wire [24:0] T_5920;
  wire [3:0] GEN_16_control_ttype;
  wire  GEN_16_control_dmode;
  wire [5:0] GEN_16_control_maskmax;
  wire [39:0] GEN_16_control_reserved;
  wire  GEN_16_control_action;
  wire  GEN_16_control_chain;
  wire [1:0] GEN_16_control_zero;
  wire [1:0] GEN_16_control_tmatch;
  wire  GEN_16_control_m;
  wire  GEN_16_control_h;
  wire  GEN_16_control_s;
  wire  GEN_16_control_u;
  wire  GEN_16_control_x;
  wire  GEN_16_control_w;
  wire  GEN_16_control_r;
  wire [38:0] GEN_16_address;
  wire [63:0] T_5921;
  wire  T_5926;
  wire [23:0] T_5930;
  wire [63:0] T_5931;
  wire  T_5932;
  wire [23:0] T_5936;
  wire [63:0] T_5937;
  wire [2:0] T_5938;
  wire [1:0] T_5939;
  wire [4:0] T_5940;
  wire [3:0] T_5941;
  wire [1:0] T_5942;
  wire [5:0] T_5943;
  wire [10:0] T_5944;
  wire [1:0] T_5945;
  wire [1:0] T_5946;
  wire [3:0] T_5947;
  wire [12:0] T_5948;
  wire [2:0] T_5949;
  wire [3:0] T_5950;
  wire [16:0] T_5951;
  wire [20:0] T_5952;
  wire [31:0] T_5953;
  wire  T_5958;
  wire  T_5960;
  wire  T_5962;
  wire  T_5964;
  wire  T_5966;
  wire  T_5968;
  wire  T_5970;
  wire  T_5972;
  wire  T_5974;
  wire  T_5976;
  wire  T_5978;
  wire  T_5980;
  wire  T_5982;
  wire  T_5984;
  wire  T_5986;
  wire  T_5988;
  wire  T_5990;
  wire  T_5992;
  wire  T_5994;
  wire  T_5996;
  wire  T_5998;
  wire  T_6000;
  wire  T_6002;
  wire  T_6004;
  wire  T_6006;
  wire  T_6008;
  wire  T_6010;
  wire  T_6012;
  wire  T_6014;
  wire  T_6016;
  wire  T_6018;
  wire  T_6020;
  wire  T_6022;
  wire  T_6024;
  wire  T_6026;
  wire  T_6028;
  wire  T_6030;
  wire  T_6032;
  wire  T_6034;
  wire  T_6036;
  wire  T_6038;
  wire  T_6040;
  wire  T_6042;
  wire  T_6044;
  wire  T_6046;
  wire  T_6048;
  wire  T_6050;
  wire  T_6052;
  wire  T_6054;
  wire  T_6056;
  wire  T_6058;
  wire  T_6060;
  wire  T_6062;
  wire  T_6064;
  wire  T_6066;
  wire  T_6068;
  wire  T_6070;
  wire  T_6072;
  wire  T_6074;
  wire  T_6076;
  wire  T_6078;
  wire  T_6080;
  wire  T_6082;
  wire  T_6084;
  wire  T_6086;
  wire  T_6088;
  wire  T_6090;
  wire  T_6092;
  wire  T_6094;
  wire  T_6096;
  wire  T_6098;
  wire  T_6100;
  wire  T_6102;
  wire  T_6104;
  wire  T_6106;
  wire  T_6108;
  wire  T_6110;
  wire  T_6112;
  wire  T_6114;
  wire  T_6116;
  wire  T_6118;
  wire  T_6119;
  wire  T_6120;
  wire  T_6121;
  wire  T_6122;
  wire  T_6123;
  wire  T_6124;
  wire  T_6125;
  wire  T_6126;
  wire  T_6127;
  wire  T_6128;
  wire  T_6129;
  wire  T_6130;
  wire  T_6131;
  wire  T_6132;
  wire  T_6133;
  wire  T_6134;
  wire  T_6135;
  wire  T_6136;
  wire  T_6137;
  wire  T_6138;
  wire  T_6139;
  wire  T_6140;
  wire  T_6141;
  wire  T_6142;
  wire  T_6143;
  wire  T_6144;
  wire  T_6145;
  wire  T_6146;
  wire  T_6147;
  wire  T_6148;
  wire  T_6149;
  wire  T_6150;
  wire  T_6151;
  wire  T_6152;
  wire  T_6153;
  wire  T_6154;
  wire  T_6155;
  wire  T_6156;
  wire  T_6157;
  wire  T_6158;
  wire  T_6159;
  wire  T_6160;
  wire  T_6161;
  wire  T_6162;
  wire  T_6163;
  wire  T_6164;
  wire  T_6165;
  wire  T_6166;
  wire  T_6167;
  wire  T_6168;
  wire  T_6169;
  wire  T_6170;
  wire  T_6171;
  wire  T_6172;
  wire  T_6173;
  wire  T_6174;
  wire  T_6175;
  wire  T_6176;
  wire  T_6177;
  wire  T_6178;
  wire  T_6179;
  wire  T_6180;
  wire  T_6181;
  wire  T_6182;
  wire  T_6183;
  wire  T_6184;
  wire  T_6185;
  wire  T_6186;
  wire  T_6187;
  wire  T_6188;
  wire  T_6189;
  wire  T_6190;
  wire  T_6191;
  wire  T_6192;
  wire  T_6193;
  wire  T_6194;
  wire  T_6195;
  wire  T_6196;
  wire  T_6197;
  wire  addr_valid;
  wire [1:0] csr_addr_priv;
  wire [11:0] T_6216;
  wire  T_6218;
  wire  T_6220;
  wire  T_6221;
  wire  T_6222;
  wire  priv_sufficient;
  wire [1:0] T_6223;
  wire [1:0] T_6224;
  wire  read_only;
  wire  T_6226;
  wire  T_6228;
  wire  wen;
  wire  T_6229;
  wire  T_6230;
  wire  T_6231;
  wire [63:0] T_6233;
  wire  T_6234;
  wire [63:0] T_6236;
  wire [63:0] T_6237;
  wire [63:0] T_6240;
  wire [63:0] T_6241;
  wire [63:0] wdata;
  wire  do_system_insn;
  wire [2:0] T_6243;
  wire [7:0] opcode;
  wire  T_6244;
  wire  insn_call;
  wire  T_6245;
  wire  insn_break;
  wire  T_6246;
  wire  insn_ret;
  wire  T_6247;
  wire  insn_sfence_vm;
  wire  T_6248;
  wire  insn_wfi;
  wire  T_6249;
  wire  T_6251;
  wire  T_6253;
  wire  T_6254;
  wire  T_6265;
  wire  T_6266;
  wire  T_6269;
  wire  T_6270;
  wire  T_6271;
  wire  T_6272;
  wire  GEN_314;
  wire  T_6275;
  wire  GEN_315;
  wire  T_6278;
  wire [3:0] GEN_3;
  wire [4:0] T_6280;
  wire [3:0] T_6281;
  wire [1:0] T_6284;
  wire [3:0] T_6285;
  wire [63:0] cause;
  wire [5:0] cause_lsbs;
  wire  T_6286;
  wire  T_6288;
  wire  causeIsDebugInt;
  wire  T_6291;
  wire  causeIsDebugTrigger;
  wire  T_6297;
  wire [1:0] T_6298;
  wire [1:0] T_6299;
  wire [3:0] T_6300;
  wire [3:0] T_6301;
  wire  T_6302;
  wire  causeIsDebugBreak;
  wire  T_6304;
  wire  T_6305;
  wire  T_6306;
  wire  T_6307;
  wire [11:0] debugTVec;
  wire [39:0] T_6322;
  wire [39:0] tvec;
  wire [39:0] epc;
  wire [39:0] T_6329;
  wire  T_6332;
  wire [1:0] T_6333;
  wire  T_6335;
  wire [1:0] T_6336;
  wire  T_6338;
  wire  T_6339;
  wire [39:0] T_6340;
  wire [39:0] T_6342;
  wire [39:0] T_6343;
  wire [63:0] T_6344;
  wire  T_6345;
  wire  T_6353;
  wire  T_6354;
  wire  T_6355;
  wire  T_6356;
  wire  T_6357;
  wire  T_6358;
  wire  T_6359;
  wire  T_6360;
  wire  T_6361;
  wire  T_6362;
  wire  T_6363;
  wire  T_6364;
  wire  T_6365;
  wire [1:0] T_6371;
  wire [1:0] T_6372;
  wire [2:0] T_6373;
  wire  GEN_316;
  wire [39:0] GEN_317;
  wire [2:0] GEN_318;
  wire [1:0] GEN_319;
  wire  T_6376;
  wire [1:0] GEN_325;
  wire [39:0] GEN_328;
  wire [39:0] GEN_329;
  wire [63:0] GEN_330;
  wire [39:0] GEN_331;
  wire  GEN_332;
  wire [1:0] GEN_333;
  wire  GEN_334;
  wire [1:0] GEN_335;
  wire  GEN_336;
  wire [39:0] GEN_337;
  wire [2:0] GEN_338;
  wire [1:0] GEN_339;
  wire [1:0] GEN_344;
  wire [1:0] GEN_346;
  wire [39:0] GEN_347;
  wire [63:0] GEN_348;
  wire [39:0] GEN_349;
  wire  GEN_350;
  wire [1:0] GEN_351;
  wire  GEN_352;
  wire [1:0] GEN_358;
  wire  GEN_359;
  wire  T_6405;
  wire  GEN_360;
  wire  GEN_362;
  wire  GEN_364;
  wire [1:0] GEN_365;
  wire [1:0] GEN_366;
  wire [1:0] GEN_370;
  wire  GEN_371;
  wire  GEN_372;
  wire  GEN_373;
  wire [1:0] GEN_374;
  wire [1:0] T_6415;
  wire [1:0] GEN_4;
  wire [2:0] T_6416;
  wire  T_6418;
  wire  T_6419;
  wire  T_6421;
  wire  T_6423;
  wire [63:0] T_6425;
  wire [63:0] T_6427;
  wire [63:0] T_6435;
  wire [63:0] T_6437;
  wire [63:0] T_6439;
  wire [63:0] T_6441;
  wire [31:0] T_6443;
  wire [12:0] T_6445;
  wire [63:0] T_6447;
  wire [63:0] T_6449;
  wire [63:0] T_6451;
  wire [63:0] T_6453;
  wire [63:0] T_6455;
  wire [63:0] T_6457;
  wire [63:0] T_6459;
  wire  T_6461;
  wire [31:0] T_6463;
  wire [39:0] T_6465;
  wire [63:0] T_6467;
  wire [63:0] GEN_5;
  wire [63:0] T_6585;
  wire [63:0] T_6586;
  wire [63:0] T_6590;
  wire [63:0] T_6591;
  wire [63:0] T_6592;
  wire [63:0] T_6593;
  wire [63:0] GEN_6;
  wire [63:0] T_6594;
  wire [63:0] GEN_7;
  wire [63:0] T_6595;
  wire [63:0] T_6596;
  wire [63:0] T_6597;
  wire [63:0] T_6598;
  wire [63:0] T_6599;
  wire [63:0] T_6600;
  wire [63:0] T_6601;
  wire [63:0] T_6602;
  wire [63:0] GEN_8;
  wire [63:0] T_6603;
  wire [63:0] GEN_9;
  wire [63:0] T_6604;
  wire [63:0] GEN_10;
  wire [63:0] T_6605;
  wire [63:0] T_6606;
  wire [63:0] T_6665;
  wire [4:0] T_6666;
  wire [4:0] GEN_375;
  wire  T_6717_debug;
  wire [1:0] T_6717_prv;
  wire  T_6717_sd;
  wire [30:0] T_6717_zero3;
  wire  T_6717_sd_rv32;
  wire [1:0] T_6717_zero2;
  wire [4:0] T_6717_vm;
  wire [3:0] T_6717_zero1;
  wire  T_6717_mxr;
  wire  T_6717_pum;
  wire  T_6717_mprv;
  wire [1:0] T_6717_xs;
  wire [1:0] T_6717_fs;
  wire [1:0] T_6717_mpp;
  wire [1:0] T_6717_hpp;
  wire  T_6717_spp;
  wire  T_6717_mpie;
  wire  T_6717_hpie;
  wire  T_6717_spie;
  wire  T_6717_upie;
  wire  T_6717_mie;
  wire  T_6717_hie;
  wire  T_6717_sie;
  wire  T_6717_uie;
  wire [66:0] T_6743;
  wire  T_6744;
  wire  T_6745;
  wire  T_6746;
  wire  T_6747;
  wire  T_6748;
  wire  T_6749;
  wire  T_6750;
  wire  T_6751;
  wire  T_6752;
  wire [1:0] T_6753;
  wire [1:0] T_6754;
  wire [1:0] T_6755;
  wire [1:0] T_6756;
  wire  T_6757;
  wire  T_6758;
  wire  T_6759;
  wire [3:0] T_6760;
  wire [4:0] T_6761;
  wire [1:0] T_6762;
  wire  T_6763;
  wire [30:0] T_6764;
  wire  T_6765;
  wire [1:0] T_6766;
  wire  T_6767;
  wire  GEN_401;
  wire  GEN_402;
  wire  T_6796_rocc;
  wire  T_6796_meip;
  wire  T_6796_heip;
  wire  T_6796_seip;
  wire  T_6796_ueip;
  wire  T_6796_mtip;
  wire  T_6796_htip;
  wire  T_6796_stip;
  wire  T_6796_utip;
  wire  T_6796_msip;
  wire  T_6796_hsip;
  wire  T_6796_ssip;
  wire  T_6796_usip;
  wire  T_6810;
  wire  T_6811;
  wire  T_6812;
  wire  T_6813;
  wire  T_6814;
  wire  T_6815;
  wire  T_6816;
  wire  T_6817;
  wire  T_6818;
  wire  T_6819;
  wire  T_6820;
  wire  T_6821;
  wire  T_6822;
  wire [63:0] GEN_11;
  wire [63:0] T_6823;
  wire [63:0] GEN_416;
  wire [63:0] T_6824;
  wire [63:0] T_6826;
  wire [63:0] T_6827;
  wire [63:0] GEN_417;
  wire [63:0] GEN_418;
  wire [61:0] T_6828;
  wire [63:0] GEN_12;
  wire [63:0] T_6829;
  wire [63:0] GEN_419;
  wire [63:0] T_6831;
  wire [63:0] GEN_420;
  wire [39:0] T_6832;
  wire [39:0] GEN_421;
  wire [57:0] T_6833;
  wire [63:0] GEN_422;
  wire [57:0] GEN_423;
  wire [63:0] GEN_424;
  wire [57:0] GEN_425;
  wire [1:0] T_6871_xdebugver;
  wire  T_6871_ndreset;
  wire  T_6871_fullreset;
  wire [11:0] T_6871_zero3;
  wire  T_6871_ebreakm;
  wire  T_6871_ebreakh;
  wire  T_6871_ebreaks;
  wire  T_6871_ebreaku;
  wire  T_6871_zero2;
  wire  T_6871_stopcycle;
  wire  T_6871_stoptime;
  wire [2:0] T_6871_cause;
  wire  T_6871_debugint;
  wire  T_6871_zero1;
  wire  T_6871_halt;
  wire  T_6871_step;
  wire [1:0] T_6871_prv;
  wire [1:0] T_6889;
  wire [2:0] T_6894;
  wire  T_6899;
  wire  T_6900;
  wire  T_6901;
  wire [11:0] T_6902;
  wire  T_6903;
  wire  T_6904;
  wire [1:0] T_6905;
  wire  GEN_443;
  wire  GEN_444;
  wire  GEN_445;
  wire [63:0] GEN_446;
  wire [63:0] GEN_447;
  wire [3:0] GEN_17_control_ttype;
  wire  GEN_17_control_dmode;
  wire [5:0] GEN_17_control_maskmax;
  wire [39:0] GEN_17_control_reserved;
  wire  GEN_17_control_action;
  wire  GEN_17_control_chain;
  wire [1:0] GEN_17_control_zero;
  wire [1:0] GEN_17_control_tmatch;
  wire  GEN_17_control_m;
  wire  GEN_17_control_h;
  wire  GEN_17_control_s;
  wire  GEN_17_control_u;
  wire  GEN_17_control_x;
  wire  GEN_17_control_w;
  wire  GEN_17_control_r;
  wire [38:0] GEN_17_address;
  wire  T_6928;
  wire  T_6929;
  wire [3:0] T_6962_ttype;
  wire  T_6962_dmode;
  wire [5:0] T_6962_maskmax;
  wire [39:0] T_6962_reserved;
  wire  T_6962_action;
  wire  T_6962_chain;
  wire [1:0] T_6962_zero;
  wire [1:0] T_6962_tmatch;
  wire  T_6962_m;
  wire  T_6962_h;
  wire  T_6962_s;
  wire  T_6962_u;
  wire  T_6962_x;
  wire  T_6962_w;
  wire  T_6962_r;
  wire [1:0] T_6985;
  wire [1:0] T_6986;
  wire [39:0] T_6989;
  wire [5:0] T_6990;
  wire  T_6991;
  wire [3:0] T_6992;
  wire  T_6993;
  wire [3:0] GEN_18;
  wire  GEN_19;
  wire  GEN_467;
  wire [5:0] GEN_20;
  wire [39:0] GEN_21;
  wire  GEN_22;
  wire  GEN_473;
  wire  GEN_23;
  wire [1:0] GEN_24;
  wire [1:0] GEN_25;
  wire [1:0] GEN_479;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_489;
  wire  GEN_31;
  wire  GEN_491;
  wire  GEN_32;
  wire  GEN_493;
  wire  GEN_33;
  wire  GEN_495;
  wire  T_6994;
  wire  GEN_34;
  wire  GEN_497;
  wire  GEN_518;
  wire  GEN_527;
  wire [1:0] GEN_536;
  wire  GEN_551;
  wire  GEN_554;
  wire  GEN_557;
  wire [38:0] GEN_35;
  wire [38:0] GEN_561;
  wire [38:0] GEN_564;
  wire  GEN_585;
  wire  GEN_594;
  wire [1:0] GEN_603;
  wire  GEN_618;
  wire  GEN_621;
  wire  GEN_624;
  wire [38:0] GEN_629;
  wire  GEN_656;
  wire  GEN_657;
  wire [63:0] GEN_671;
  wire [63:0] GEN_672;
  wire [63:0] GEN_673;
  wire [63:0] GEN_674;
  wire [63:0] GEN_675;
  wire [39:0] GEN_676;
  wire [63:0] GEN_677;
  wire [57:0] GEN_678;
  wire [63:0] GEN_679;
  wire [57:0] GEN_680;
  wire  GEN_698;
  wire  GEN_699;
  wire  GEN_700;
  wire [63:0] GEN_701;
  wire [63:0] GEN_702;
  wire  GEN_739;
  wire  GEN_748;
  wire [1:0] GEN_757;
  wire  GEN_772;
  wire  GEN_775;
  wire  GEN_778;
  wire [38:0] GEN_783;
  wire  GEN_785;
  wire  GEN_786;
  wire  GEN_787;
  wire  GEN_788;
  wire  GEN_789;
  wire [3:0] T_7061_control_ttype;
  wire  T_7061_control_dmode;
  wire [5:0] T_7061_control_maskmax;
  wire [39:0] T_7061_control_reserved;
  wire  T_7061_control_action;
  wire  T_7061_control_chain;
  wire [1:0] T_7061_control_zero;
  wire [1:0] T_7061_control_tmatch;
  wire  T_7061_control_m;
  wire  T_7061_control_h;
  wire  T_7061_control_s;
  wire  T_7061_control_u;
  wire  T_7061_control_x;
  wire  T_7061_control_w;
  wire  T_7061_control_r;
  wire [38:0] T_7061_address;
  wire [102:0] T_7080;
  wire [38:0] T_7081;
  wire  T_7082;
  wire  T_7083;
  wire  T_7084;
  wire  T_7085;
  wire  T_7086;
  wire  T_7087;
  wire  T_7088;
  wire [1:0] T_7089;
  wire [1:0] T_7090;
  wire  T_7091;
  wire  T_7092;
  wire [39:0] T_7093;
  wire [5:0] T_7094;
  wire  T_7095;
  wire [3:0] T_7096;
  wire  GEN_13;
  reg [31:0] GEN_235;
  wire [6:0] GEN_14;
  reg [31:0] GEN_236;
  wire [4:0] GEN_15;
  reg [31:0] GEN_237;
  wire [4:0] GEN_16;
  reg [31:0] GEN_238;
  wire  GEN_17;
  reg [31:0] GEN_239;
  wire  GEN_58;
  reg [31:0] GEN_240;
  wire  GEN_59;
  reg [31:0] GEN_241;
  wire [4:0] GEN_60;
  reg [31:0] GEN_242;
  wire [6:0] GEN_61;
  reg [31:0] GEN_243;
  wire [63:0] GEN_62;
  reg [63:0] GEN_244;
  wire [63:0] GEN_63;
  reg [63:0] GEN_245;
  wire  GEN_64;
  reg [31:0] GEN_246;
  wire [1:0] GEN_65;
  reg [31:0] GEN_247;
  wire  GEN_66;
  reg [31:0] GEN_248;
  wire [30:0] GEN_67;
  reg [31:0] GEN_249;
  wire  GEN_68;
  reg [31:0] GEN_250;
  wire [1:0] GEN_69;
  reg [31:0] GEN_251;
  wire [4:0] GEN_70;
  reg [31:0] GEN_252;
  wire [3:0] GEN_71;
  reg [31:0] GEN_253;
  wire  GEN_72;
  reg [31:0] GEN_254;
  wire  GEN_73;
  reg [31:0] GEN_255;
  wire  GEN_74;
  reg [31:0] GEN_256;
  wire [1:0] GEN_75;
  reg [31:0] GEN_257;
  wire [1:0] GEN_76;
  reg [31:0] GEN_258;
  wire [1:0] GEN_77;
  reg [31:0] GEN_259;
  wire [1:0] GEN_78;
  reg [31:0] GEN_260;
  wire  GEN_79;
  reg [31:0] GEN_261;
  wire  GEN_80;
  reg [31:0] GEN_262;
  wire  GEN_81;
  reg [31:0] GEN_263;
  wire  GEN_82;
  reg [31:0] GEN_264;
  wire  GEN_83;
  reg [31:0] GEN_265;
  wire  GEN_84;
  reg [31:0] GEN_266;
  wire  GEN_85;
  reg [31:0] GEN_267;
  wire  GEN_86;
  reg [31:0] GEN_268;
  wire  GEN_87;
  reg [31:0] GEN_269;
  wire  GEN_88;
  reg [31:0] GEN_270;
  wire  GEN_89;
  reg [31:0] GEN_271;
  wire  GEN_90;
  reg [31:0] GEN_272;
  wire  GEN_91;
  reg [31:0] GEN_273;
  wire [39:0] GEN_92;
  reg [63:0] GEN_274;
  wire [5:0] GEN_93;
  reg [31:0] GEN_275;
  wire [4:0] GEN_94;
  reg [31:0] GEN_276;
  wire [2:0] GEN_95;
  reg [31:0] GEN_277;
  wire [63:0] GEN_96;
  reg [63:0] GEN_278;
  wire  GEN_97;
  reg [31:0] GEN_279;
  wire  GEN_98;
  reg [31:0] GEN_280;
  wire [63:0] GEN_99;
  reg [63:0] GEN_281;
  wire [63:0] GEN_100;
  reg [63:0] GEN_282;
  wire  GEN_101;
  reg [31:0] GEN_283;
  wire  GEN_102;
  reg [31:0] GEN_284;
  wire  GEN_103;
  reg [31:0] GEN_285;
  wire  GEN_104;
  reg [31:0] GEN_286;
  wire  GEN_105;
  reg [31:0] GEN_287;
  wire  GEN_106;
  reg [31:0] GEN_288;
  wire  GEN_107;
  reg [31:0] GEN_289;
  wire  GEN_108;
  reg [31:0] GEN_290;
  wire [2:0] GEN_109;
  reg [31:0] GEN_291;
  wire  GEN_110;
  reg [31:0] GEN_292;
  wire [1:0] GEN_111;
  reg [31:0] GEN_293;
  wire  GEN_112;
  reg [31:0] GEN_294;
  wire [3:0] GEN_113;
  reg [31:0] GEN_295;
  wire [63:0] GEN_114;
  reg [63:0] GEN_296;
  wire  GEN_115;
  reg [31:0] GEN_297;
  wire  GEN_116;
  reg [31:0] GEN_298;
  wire [64:0] GEN_117;
  reg [95:0] GEN_299;
  wire [4:0] GEN_118;
  reg [31:0] GEN_300;
  wire  GEN_119;
  reg [31:0] GEN_301;
  assign io_rw_rdata = T_6665;
  assign io_csr_stall = reg_wfi;
  assign io_csr_xcpt = T_6272;
  assign io_eret = insn_ret;
  assign io_singleStep = T_6332;
  assign io_status_debug = reg_debug;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_sd = T_6339;
  assign io_status_zero3 = reg_mstatus_zero3;
  assign io_status_sd_rv32 = reg_mstatus_sd_rv32;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign io_status_vm = reg_mstatus_vm;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign io_status_mxr = reg_mstatus_mxr;
  assign io_status_pum = reg_mstatus_pum;
  assign io_status_mprv = reg_mstatus_mprv;
  assign io_status_xs = reg_mstatus_xs;
  assign io_status_fs = reg_mstatus_fs;
  assign io_status_mpp = reg_mstatus_mpp;
  assign io_status_hpp = reg_mstatus_hpp;
  assign io_status_spp = reg_mstatus_spp;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_hpie = reg_mstatus_hpie;
  assign io_status_spie = reg_mstatus_spie;
  assign io_status_upie = reg_mstatus_upie;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_hie = reg_mstatus_hie;
  assign io_status_sie = reg_mstatus_sie;
  assign io_status_uie = reg_mstatus_uie;
  assign io_ptbr_asid = reg_sptbr_asid;
  assign io_ptbr_ppn = reg_sptbr_ppn;
  assign io_evec = T_6329;
  assign io_fatc = insn_sfence_vm;
  assign io_time = T_5586;
  assign io_fcsr_rm = reg_frm;
  assign io_rocc_cmd_valid = GEN_13;
  assign io_rocc_cmd_bits_inst_funct = GEN_14;
  assign io_rocc_cmd_bits_inst_rs2 = GEN_15;
  assign io_rocc_cmd_bits_inst_rs1 = GEN_16;
  assign io_rocc_cmd_bits_inst_xd = GEN_17;
  assign io_rocc_cmd_bits_inst_xs1 = GEN_58;
  assign io_rocc_cmd_bits_inst_xs2 = GEN_59;
  assign io_rocc_cmd_bits_inst_rd = GEN_60;
  assign io_rocc_cmd_bits_inst_opcode = GEN_61;
  assign io_rocc_cmd_bits_rs1 = GEN_62;
  assign io_rocc_cmd_bits_rs2 = GEN_63;
  assign io_rocc_cmd_bits_status_debug = GEN_64;
  assign io_rocc_cmd_bits_status_prv = GEN_65;
  assign io_rocc_cmd_bits_status_sd = GEN_66;
  assign io_rocc_cmd_bits_status_zero3 = GEN_67;
  assign io_rocc_cmd_bits_status_sd_rv32 = GEN_68;
  assign io_rocc_cmd_bits_status_zero2 = GEN_69;
  assign io_rocc_cmd_bits_status_vm = GEN_70;
  assign io_rocc_cmd_bits_status_zero1 = GEN_71;
  assign io_rocc_cmd_bits_status_mxr = GEN_72;
  assign io_rocc_cmd_bits_status_pum = GEN_73;
  assign io_rocc_cmd_bits_status_mprv = GEN_74;
  assign io_rocc_cmd_bits_status_xs = GEN_75;
  assign io_rocc_cmd_bits_status_fs = GEN_76;
  assign io_rocc_cmd_bits_status_mpp = GEN_77;
  assign io_rocc_cmd_bits_status_hpp = GEN_78;
  assign io_rocc_cmd_bits_status_spp = GEN_79;
  assign io_rocc_cmd_bits_status_mpie = GEN_80;
  assign io_rocc_cmd_bits_status_hpie = GEN_81;
  assign io_rocc_cmd_bits_status_spie = GEN_82;
  assign io_rocc_cmd_bits_status_upie = GEN_83;
  assign io_rocc_cmd_bits_status_mie = GEN_84;
  assign io_rocc_cmd_bits_status_hie = GEN_85;
  assign io_rocc_cmd_bits_status_sie = GEN_86;
  assign io_rocc_cmd_bits_status_uie = GEN_87;
  assign io_rocc_resp_ready = GEN_88;
  assign io_rocc_mem_req_ready = GEN_89;
  assign io_rocc_mem_s2_nack = GEN_90;
  assign io_rocc_mem_resp_valid = GEN_91;
  assign io_rocc_mem_resp_bits_addr = GEN_92;
  assign io_rocc_mem_resp_bits_tag = GEN_93;
  assign io_rocc_mem_resp_bits_cmd = GEN_94;
  assign io_rocc_mem_resp_bits_typ = GEN_95;
  assign io_rocc_mem_resp_bits_data = GEN_96;
  assign io_rocc_mem_resp_bits_replay = GEN_97;
  assign io_rocc_mem_resp_bits_has_data = GEN_98;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_99;
  assign io_rocc_mem_resp_bits_store_data = GEN_100;
  assign io_rocc_mem_replay_next = GEN_101;
  assign io_rocc_mem_xcpt_ma_ld = GEN_102;
  assign io_rocc_mem_xcpt_ma_st = GEN_103;
  assign io_rocc_mem_xcpt_pf_ld = GEN_104;
  assign io_rocc_mem_xcpt_pf_st = GEN_105;
  assign io_rocc_mem_ordered = GEN_106;
  assign io_rocc_autl_acquire_ready = GEN_107;
  assign io_rocc_autl_grant_valid = GEN_108;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_109;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_110;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_111;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_112;
  assign io_rocc_autl_grant_bits_g_type = GEN_113;
  assign io_rocc_autl_grant_bits_data = GEN_114;
  assign io_rocc_fpu_req_ready = GEN_115;
  assign io_rocc_fpu_resp_valid = GEN_116;
  assign io_rocc_fpu_resp_bits_data = GEN_117;
  assign io_rocc_fpu_resp_bits_exc = GEN_118;
  assign io_rocc_exception = GEN_119;
  assign io_interrupt = GEN_40;
  assign io_interrupt_cause = GEN_41;
  assign io_bp_0_control_ttype = reg_bp_0_control_ttype;
  assign io_bp_0_control_dmode = reg_bp_0_control_dmode;
  assign io_bp_0_control_maskmax = reg_bp_0_control_maskmax;
  assign io_bp_0_control_reserved = reg_bp_0_control_reserved;
  assign io_bp_0_control_action = reg_bp_0_control_action;
  assign io_bp_0_control_chain = reg_bp_0_control_chain;
  assign io_bp_0_control_zero = reg_bp_0_control_zero;
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch;
  assign io_bp_0_control_m = reg_bp_0_control_m;
  assign io_bp_0_control_h = reg_bp_0_control_h;
  assign io_bp_0_control_s = reg_bp_0_control_s;
  assign io_bp_0_control_u = reg_bp_0_control_u;
  assign io_bp_0_control_x = reg_bp_0_control_x;
  assign io_bp_0_control_w = reg_bp_0_control_w;
  assign io_bp_0_control_r = reg_bp_0_control_r;
  assign io_bp_0_address = reg_bp_0_address;
  assign T_4982_debug = T_5032;
  assign T_4982_prv = T_5031;
  assign T_4982_sd = T_5030;
  assign T_4982_zero3 = T_5029;
  assign T_4982_sd_rv32 = T_5028;
  assign T_4982_zero2 = T_5027;
  assign T_4982_vm = T_5026;
  assign T_4982_zero1 = T_5025;
  assign T_4982_mxr = T_5024;
  assign T_4982_pum = T_5023;
  assign T_4982_mprv = T_5022;
  assign T_4982_xs = T_5021;
  assign T_4982_fs = T_5020;
  assign T_4982_mpp = T_5019;
  assign T_4982_hpp = T_5018;
  assign T_4982_spp = T_5017;
  assign T_4982_mpie = T_5016;
  assign T_4982_hpie = T_5015;
  assign T_4982_spie = T_5014;
  assign T_4982_upie = T_5013;
  assign T_4982_mie = T_5012;
  assign T_4982_hie = T_5011;
  assign T_4982_sie = T_5010;
  assign T_4982_uie = T_5009;
  assign T_5008 = 67'h0;
  assign T_5009 = T_5008[0];
  assign T_5010 = T_5008[1];
  assign T_5011 = T_5008[2];
  assign T_5012 = T_5008[3];
  assign T_5013 = T_5008[4];
  assign T_5014 = T_5008[5];
  assign T_5015 = T_5008[6];
  assign T_5016 = T_5008[7];
  assign T_5017 = T_5008[8];
  assign T_5018 = T_5008[10:9];
  assign T_5019 = T_5008[12:11];
  assign T_5020 = T_5008[14:13];
  assign T_5021 = T_5008[16:15];
  assign T_5022 = T_5008[17];
  assign T_5023 = T_5008[18];
  assign T_5024 = T_5008[19];
  assign T_5025 = T_5008[23:20];
  assign T_5026 = T_5008[28:24];
  assign T_5027 = T_5008[30:29];
  assign T_5028 = T_5008[31];
  assign T_5029 = T_5008[62:32];
  assign T_5030 = T_5008[63];
  assign T_5031 = T_5008[65:64];
  assign T_5032 = T_5008[66];
  assign reset_mstatus_debug = T_4982_debug;
  assign reset_mstatus_prv = 2'h3;
  assign reset_mstatus_sd = T_4982_sd;
  assign reset_mstatus_zero3 = T_4982_zero3;
  assign reset_mstatus_sd_rv32 = T_4982_sd_rv32;
  assign reset_mstatus_zero2 = T_4982_zero2;
  assign reset_mstatus_vm = T_4982_vm;
  assign reset_mstatus_zero1 = T_4982_zero1;
  assign reset_mstatus_mxr = T_4982_mxr;
  assign reset_mstatus_pum = T_4982_pum;
  assign reset_mstatus_mprv = T_4982_mprv;
  assign reset_mstatus_xs = T_4982_xs;
  assign reset_mstatus_fs = T_4982_fs;
  assign reset_mstatus_mpp = 2'h3;
  assign reset_mstatus_hpp = T_4982_hpp;
  assign reset_mstatus_spp = T_4982_spp;
  assign reset_mstatus_mpie = T_4982_mpie;
  assign reset_mstatus_hpie = T_4982_hpie;
  assign reset_mstatus_spie = T_4982_spie;
  assign reset_mstatus_upie = T_4982_upie;
  assign reset_mstatus_mie = T_4982_mie;
  assign reset_mstatus_hie = T_4982_hie;
  assign reset_mstatus_sie = T_4982_sie;
  assign reset_mstatus_uie = T_4982_uie;
  assign new_prv = GEN_370;
  assign T_5121_xdebugver = T_5157;
  assign T_5121_ndreset = T_5156;
  assign T_5121_fullreset = T_5155;
  assign T_5121_zero3 = T_5154;
  assign T_5121_ebreakm = T_5153;
  assign T_5121_ebreakh = T_5152;
  assign T_5121_ebreaks = T_5151;
  assign T_5121_ebreaku = T_5150;
  assign T_5121_zero2 = T_5149;
  assign T_5121_stopcycle = T_5148;
  assign T_5121_stoptime = T_5147;
  assign T_5121_cause = T_5146;
  assign T_5121_debugint = T_5145;
  assign T_5121_zero1 = T_5144;
  assign T_5121_halt = T_5143;
  assign T_5121_step = T_5142;
  assign T_5121_prv = T_5141;
  assign T_5140 = 32'h0;
  assign T_5141 = T_5140[1:0];
  assign T_5142 = T_5140[2];
  assign T_5143 = T_5140[3];
  assign T_5144 = T_5140[4];
  assign T_5145 = T_5140[5];
  assign T_5146 = T_5140[8:6];
  assign T_5147 = T_5140[9];
  assign T_5148 = T_5140[10];
  assign T_5149 = T_5140[11];
  assign T_5150 = T_5140[12];
  assign T_5151 = T_5140[13];
  assign T_5152 = T_5140[14];
  assign T_5153 = T_5140[15];
  assign T_5154 = T_5140[27:16];
  assign T_5155 = T_5140[28];
  assign T_5156 = T_5140[29];
  assign T_5157 = T_5140[31:30];
  assign reset_dcsr_xdebugver = 2'h1;
  assign reset_dcsr_ndreset = T_5121_ndreset;
  assign reset_dcsr_fullreset = T_5121_fullreset;
  assign reset_dcsr_zero3 = T_5121_zero3;
  assign reset_dcsr_ebreakm = T_5121_ebreakm;
  assign reset_dcsr_ebreakh = T_5121_ebreakh;
  assign reset_dcsr_ebreaks = T_5121_ebreaks;
  assign reset_dcsr_ebreaku = T_5121_ebreaku;
  assign reset_dcsr_zero2 = T_5121_zero2;
  assign reset_dcsr_stopcycle = T_5121_stopcycle;
  assign reset_dcsr_stoptime = T_5121_stoptime;
  assign reset_dcsr_cause = T_5121_cause;
  assign reset_dcsr_debugint = T_5121_debugint;
  assign reset_dcsr_zero1 = T_5121_zero1;
  assign reset_dcsr_halt = T_5121_halt;
  assign reset_dcsr_step = T_5121_step;
  assign reset_dcsr_prv = 2'h3;
  assign T_5223_rocc = T_5251;
  assign T_5223_meip = T_5250;
  assign T_5223_heip = T_5249;
  assign T_5223_seip = T_5248;
  assign T_5223_ueip = T_5247;
  assign T_5223_mtip = T_5246;
  assign T_5223_htip = T_5245;
  assign T_5223_stip = T_5244;
  assign T_5223_utip = T_5243;
  assign T_5223_msip = T_5242;
  assign T_5223_hsip = T_5241;
  assign T_5223_ssip = T_5240;
  assign T_5223_usip = T_5239;
  assign T_5238 = 13'h0;
  assign T_5239 = T_5238[0];
  assign T_5240 = T_5238[1];
  assign T_5241 = T_5238[2];
  assign T_5242 = T_5238[3];
  assign T_5243 = T_5238[4];
  assign T_5244 = T_5238[5];
  assign T_5245 = T_5238[6];
  assign T_5246 = T_5238[7];
  assign T_5247 = T_5238[8];
  assign T_5248 = T_5238[9];
  assign T_5249 = T_5238[10];
  assign T_5250 = T_5238[11];
  assign T_5251 = T_5238[12];
  assign T_5252_rocc = 1'h0;
  assign T_5252_meip = 1'h1;
  assign T_5252_heip = T_5223_heip;
  assign T_5252_seip = 1'h0;
  assign T_5252_ueip = T_5223_ueip;
  assign T_5252_mtip = 1'h1;
  assign T_5252_htip = T_5223_htip;
  assign T_5252_stip = 1'h0;
  assign T_5252_utip = T_5223_utip;
  assign T_5252_msip = 1'h1;
  assign T_5252_hsip = T_5223_hsip;
  assign T_5252_ssip = 1'h0;
  assign T_5252_usip = T_5223_usip;
  assign T_5273_rocc = T_5252_rocc;
  assign T_5273_meip = 1'h0;
  assign T_5273_heip = T_5252_heip;
  assign T_5273_seip = T_5252_seip;
  assign T_5273_ueip = T_5252_ueip;
  assign T_5273_mtip = 1'h0;
  assign T_5273_htip = T_5252_htip;
  assign T_5273_stip = T_5252_stip;
  assign T_5273_utip = T_5252_utip;
  assign T_5273_msip = 1'h0;
  assign T_5273_hsip = T_5252_hsip;
  assign T_5273_ssip = T_5252_ssip;
  assign T_5273_usip = T_5252_usip;
  assign T_5290 = {T_5252_hsip,T_5252_ssip};
  assign T_5291 = {T_5290,T_5252_usip};
  assign T_5292 = {T_5252_stip,T_5252_utip};
  assign T_5293 = {T_5292,T_5252_msip};
  assign T_5294 = {T_5293,T_5291};
  assign T_5295 = {T_5252_ueip,T_5252_mtip};
  assign T_5296 = {T_5295,T_5252_htip};
  assign T_5297 = {T_5252_heip,T_5252_seip};
  assign T_5298 = {T_5252_rocc,T_5252_meip};
  assign T_5299 = {T_5298,T_5297};
  assign T_5300 = {T_5299,T_5296};
  assign supported_interrupts = {T_5300,T_5294};
  assign exception = io_exception | io_csr_xcpt;
  assign T_5317 = io_retire | exception;
  assign GEN_36 = T_5317 ? 1'h1 : reg_singleStepped;
  assign T_5320 = io_singleStep == 1'h0;
  assign GEN_37 = T_5320 ? 1'h0 : GEN_36;
  assign T_5331 = reg_singleStepped == 1'h0;
  assign T_5333 = io_retire == 1'h0;
  assign T_5334 = T_5331 | T_5333;
  assign T_5335 = T_5334 | reset;
  assign T_5337 = T_5335 == 1'h0;
  assign GEN_0 = {{5'd0}, io_retire};
  assign T_5568 = T_5567 + GEN_0;
  assign T_5571 = T_5568[6];
  assign T_5573 = T_5570 + 58'h1;
  assign T_5574 = T_5573[57:0];
  assign GEN_38 = T_5571 ? T_5574 : T_5570;
  assign T_5575 = {T_5570,T_5567};
  assign T_5579 = T_5578 + 6'h1;
  assign T_5582 = T_5579[6];
  assign T_5584 = T_5581 + 58'h1;
  assign T_5585 = T_5584[57:0];
  assign GEN_39 = T_5582 ? T_5585 : T_5581;
  assign T_5586 = {T_5581,T_5578};
  assign mip_rocc = io_rocc_interrupt;
  assign mip_meip = reg_mip_meip;
  assign mip_heip = reg_mip_heip;
  assign mip_seip = reg_mip_seip;
  assign mip_ueip = reg_mip_ueip;
  assign mip_mtip = reg_mip_mtip;
  assign mip_htip = reg_mip_htip;
  assign mip_stip = reg_mip_stip;
  assign mip_utip = reg_mip_utip;
  assign mip_msip = reg_mip_msip;
  assign mip_hsip = reg_mip_hsip;
  assign mip_ssip = reg_mip_ssip;
  assign mip_usip = reg_mip_usip;
  assign T_5600 = {mip_hsip,mip_ssip};
  assign T_5601 = {T_5600,mip_usip};
  assign T_5602 = {mip_stip,mip_utip};
  assign T_5603 = {T_5602,mip_msip};
  assign T_5604 = {T_5603,T_5601};
  assign T_5605 = {mip_ueip,mip_mtip};
  assign T_5606 = {T_5605,mip_htip};
  assign T_5607 = {mip_heip,mip_seip};
  assign T_5608 = {mip_rocc,mip_meip};
  assign T_5609 = {T_5608,T_5607};
  assign T_5610 = {T_5609,T_5606};
  assign T_5611 = {T_5610,T_5604};
  assign read_mip = T_5611 & supported_interrupts;
  assign GEN_1 = {{51'd0}, read_mip};
  assign pending_interrupts = GEN_1 & reg_mie;
  assign T_5613 = reg_debug == 1'h0;
  assign T_5615 = reg_mstatus_prv < 2'h3;
  assign T_5617 = reg_mstatus_prv == 2'h3;
  assign T_5618 = T_5617 & reg_mstatus_mie;
  assign T_5619 = T_5615 | T_5618;
  assign T_5620 = T_5613 & T_5619;
  assign T_5621 = ~ reg_mideleg;
  assign T_5622 = pending_interrupts & T_5621;
  assign m_interrupts = T_5620 ? T_5622 : 64'h0;
  assign T_5627 = reg_mstatus_prv < 2'h1;
  assign T_5629 = reg_mstatus_prv == 2'h1;
  assign T_5630 = T_5629 & reg_mstatus_sie;
  assign T_5631 = T_5627 | T_5630;
  assign T_5632 = T_5613 & T_5631;
  assign T_5633 = pending_interrupts & reg_mideleg;
  assign s_interrupts = T_5632 ? T_5633 : 64'h0;
  assign all_interrupts = m_interrupts | s_interrupts;
  assign T_5636 = all_interrupts[0];
  assign T_5637 = all_interrupts[1];
  assign T_5638 = all_interrupts[2];
  assign T_5639 = all_interrupts[3];
  assign T_5640 = all_interrupts[4];
  assign T_5641 = all_interrupts[5];
  assign T_5642 = all_interrupts[6];
  assign T_5643 = all_interrupts[7];
  assign T_5644 = all_interrupts[8];
  assign T_5645 = all_interrupts[9];
  assign T_5646 = all_interrupts[10];
  assign T_5647 = all_interrupts[11];
  assign T_5648 = all_interrupts[12];
  assign T_5649 = all_interrupts[13];
  assign T_5650 = all_interrupts[14];
  assign T_5651 = all_interrupts[15];
  assign T_5652 = all_interrupts[16];
  assign T_5653 = all_interrupts[17];
  assign T_5654 = all_interrupts[18];
  assign T_5655 = all_interrupts[19];
  assign T_5656 = all_interrupts[20];
  assign T_5657 = all_interrupts[21];
  assign T_5658 = all_interrupts[22];
  assign T_5659 = all_interrupts[23];
  assign T_5660 = all_interrupts[24];
  assign T_5661 = all_interrupts[25];
  assign T_5662 = all_interrupts[26];
  assign T_5663 = all_interrupts[27];
  assign T_5664 = all_interrupts[28];
  assign T_5665 = all_interrupts[29];
  assign T_5666 = all_interrupts[30];
  assign T_5667 = all_interrupts[31];
  assign T_5668 = all_interrupts[32];
  assign T_5669 = all_interrupts[33];
  assign T_5670 = all_interrupts[34];
  assign T_5671 = all_interrupts[35];
  assign T_5672 = all_interrupts[36];
  assign T_5673 = all_interrupts[37];
  assign T_5674 = all_interrupts[38];
  assign T_5675 = all_interrupts[39];
  assign T_5676 = all_interrupts[40];
  assign T_5677 = all_interrupts[41];
  assign T_5678 = all_interrupts[42];
  assign T_5679 = all_interrupts[43];
  assign T_5680 = all_interrupts[44];
  assign T_5681 = all_interrupts[45];
  assign T_5682 = all_interrupts[46];
  assign T_5683 = all_interrupts[47];
  assign T_5684 = all_interrupts[48];
  assign T_5685 = all_interrupts[49];
  assign T_5686 = all_interrupts[50];
  assign T_5687 = all_interrupts[51];
  assign T_5688 = all_interrupts[52];
  assign T_5689 = all_interrupts[53];
  assign T_5690 = all_interrupts[54];
  assign T_5691 = all_interrupts[55];
  assign T_5692 = all_interrupts[56];
  assign T_5693 = all_interrupts[57];
  assign T_5694 = all_interrupts[58];
  assign T_5695 = all_interrupts[59];
  assign T_5696 = all_interrupts[60];
  assign T_5697 = all_interrupts[61];
  assign T_5698 = all_interrupts[62];
  assign T_5764 = T_5698 ? 6'h3e : 6'h3f;
  assign T_5765 = T_5697 ? 6'h3d : T_5764;
  assign T_5766 = T_5696 ? 6'h3c : T_5765;
  assign T_5767 = T_5695 ? 6'h3b : T_5766;
  assign T_5768 = T_5694 ? 6'h3a : T_5767;
  assign T_5769 = T_5693 ? 6'h39 : T_5768;
  assign T_5770 = T_5692 ? 6'h38 : T_5769;
  assign T_5771 = T_5691 ? 6'h37 : T_5770;
  assign T_5772 = T_5690 ? 6'h36 : T_5771;
  assign T_5773 = T_5689 ? 6'h35 : T_5772;
  assign T_5774 = T_5688 ? 6'h34 : T_5773;
  assign T_5775 = T_5687 ? 6'h33 : T_5774;
  assign T_5776 = T_5686 ? 6'h32 : T_5775;
  assign T_5777 = T_5685 ? 6'h31 : T_5776;
  assign T_5778 = T_5684 ? 6'h30 : T_5777;
  assign T_5779 = T_5683 ? 6'h2f : T_5778;
  assign T_5780 = T_5682 ? 6'h2e : T_5779;
  assign T_5781 = T_5681 ? 6'h2d : T_5780;
  assign T_5782 = T_5680 ? 6'h2c : T_5781;
  assign T_5783 = T_5679 ? 6'h2b : T_5782;
  assign T_5784 = T_5678 ? 6'h2a : T_5783;
  assign T_5785 = T_5677 ? 6'h29 : T_5784;
  assign T_5786 = T_5676 ? 6'h28 : T_5785;
  assign T_5787 = T_5675 ? 6'h27 : T_5786;
  assign T_5788 = T_5674 ? 6'h26 : T_5787;
  assign T_5789 = T_5673 ? 6'h25 : T_5788;
  assign T_5790 = T_5672 ? 6'h24 : T_5789;
  assign T_5791 = T_5671 ? 6'h23 : T_5790;
  assign T_5792 = T_5670 ? 6'h22 : T_5791;
  assign T_5793 = T_5669 ? 6'h21 : T_5792;
  assign T_5794 = T_5668 ? 6'h20 : T_5793;
  assign T_5795 = T_5667 ? 6'h1f : T_5794;
  assign T_5796 = T_5666 ? 6'h1e : T_5795;
  assign T_5797 = T_5665 ? 6'h1d : T_5796;
  assign T_5798 = T_5664 ? 6'h1c : T_5797;
  assign T_5799 = T_5663 ? 6'h1b : T_5798;
  assign T_5800 = T_5662 ? 6'h1a : T_5799;
  assign T_5801 = T_5661 ? 6'h19 : T_5800;
  assign T_5802 = T_5660 ? 6'h18 : T_5801;
  assign T_5803 = T_5659 ? 6'h17 : T_5802;
  assign T_5804 = T_5658 ? 6'h16 : T_5803;
  assign T_5805 = T_5657 ? 6'h15 : T_5804;
  assign T_5806 = T_5656 ? 6'h14 : T_5805;
  assign T_5807 = T_5655 ? 6'h13 : T_5806;
  assign T_5808 = T_5654 ? 6'h12 : T_5807;
  assign T_5809 = T_5653 ? 6'h11 : T_5808;
  assign T_5810 = T_5652 ? 6'h10 : T_5809;
  assign T_5811 = T_5651 ? 6'hf : T_5810;
  assign T_5812 = T_5650 ? 6'he : T_5811;
  assign T_5813 = T_5649 ? 6'hd : T_5812;
  assign T_5814 = T_5648 ? 6'hc : T_5813;
  assign T_5815 = T_5647 ? 6'hb : T_5814;
  assign T_5816 = T_5646 ? 6'ha : T_5815;
  assign T_5817 = T_5645 ? 6'h9 : T_5816;
  assign T_5818 = T_5644 ? 6'h8 : T_5817;
  assign T_5819 = T_5643 ? 6'h7 : T_5818;
  assign T_5820 = T_5642 ? 6'h6 : T_5819;
  assign T_5821 = T_5641 ? 6'h5 : T_5820;
  assign T_5822 = T_5640 ? 6'h4 : T_5821;
  assign T_5823 = T_5639 ? 6'h3 : T_5822;
  assign T_5824 = T_5638 ? 6'h2 : T_5823;
  assign T_5825 = T_5637 ? 6'h1 : T_5824;
  assign T_5826 = T_5636 ? 6'h0 : T_5825;
  assign GEN_2 = {{58'd0}, T_5826};
  assign T_5827 = 64'h8000000000000000 + GEN_2;
  assign interruptCause = T_5827[63:0];
  assign T_5829 = all_interrupts != 64'h0;
  assign T_5832 = T_5829 & T_5320;
  assign T_5833 = T_5832 | reg_singleStepped;
  assign T_5838 = reg_dcsr_debugint & T_5613;
  assign GEN_40 = T_5838 ? 1'h1 : T_5833;
  assign GEN_41 = T_5838 ? 64'h800000000000000d : interruptCause;
  assign system_insn = io_rw_cmd == 3'h4;
  assign T_5841 = io_rw_cmd != 3'h0;
  assign T_5843 = system_insn == 1'h0;
  assign cpu_ren = T_5841 & T_5843;
  assign T_5844 = io_rw_cmd != 3'h5;
  assign cpu_wen = cpu_ren & T_5844;
  assign T_5845 = {io_status_hie,io_status_sie};
  assign T_5846 = {T_5845,io_status_uie};
  assign T_5847 = {io_status_spie,io_status_upie};
  assign T_5848 = {T_5847,io_status_mie};
  assign T_5849 = {T_5848,T_5846};
  assign T_5850 = {io_status_spp,io_status_mpie};
  assign T_5851 = {T_5850,io_status_hpie};
  assign T_5852 = {io_status_fs,io_status_mpp};
  assign T_5853 = {T_5852,io_status_hpp};
  assign T_5854 = {T_5853,T_5851};
  assign T_5855 = {T_5854,T_5849};
  assign T_5856 = {io_status_pum,io_status_mprv};
  assign T_5857 = {T_5856,io_status_xs};
  assign T_5858 = {io_status_vm,io_status_zero1};
  assign T_5859 = {T_5858,io_status_mxr};
  assign T_5860 = {T_5859,T_5857};
  assign T_5861 = {io_status_zero3,io_status_sd_rv32};
  assign T_5862 = {T_5861,io_status_zero2};
  assign T_5863 = {io_status_debug,io_status_prv};
  assign T_5864 = {T_5863,io_status_sd};
  assign T_5865 = {T_5864,T_5862};
  assign T_5866 = {T_5865,T_5860};
  assign T_5867 = {T_5866,T_5855};
  assign read_mstatus = T_5867[63:0];
  assign GEN_0_control_ttype = GEN_42;
  assign GEN_0_control_dmode = GEN_43;
  assign GEN_0_control_maskmax = GEN_44;
  assign GEN_0_control_reserved = GEN_45;
  assign GEN_0_control_action = GEN_46;
  assign GEN_0_control_chain = GEN_47;
  assign GEN_0_control_zero = GEN_48;
  assign GEN_0_control_tmatch = GEN_49;
  assign GEN_0_control_m = GEN_50;
  assign GEN_0_control_h = GEN_51;
  assign GEN_0_control_s = GEN_52;
  assign GEN_0_control_u = GEN_53;
  assign GEN_0_control_x = GEN_54;
  assign GEN_0_control_w = GEN_55;
  assign GEN_0_control_r = GEN_56;
  assign GEN_0_address = GEN_57;
  assign GEN_42 = reg_tselect ? reg_bp_1_control_ttype : reg_bp_0_control_ttype;
  assign GEN_43 = reg_tselect ? reg_bp_1_control_dmode : reg_bp_0_control_dmode;
  assign GEN_44 = reg_tselect ? reg_bp_1_control_maskmax : reg_bp_0_control_maskmax;
  assign GEN_45 = reg_tselect ? reg_bp_1_control_reserved : reg_bp_0_control_reserved;
  assign GEN_46 = reg_tselect ? reg_bp_1_control_action : reg_bp_0_control_action;
  assign GEN_47 = reg_tselect ? reg_bp_1_control_chain : reg_bp_0_control_chain;
  assign GEN_48 = reg_tselect ? reg_bp_1_control_zero : reg_bp_0_control_zero;
  assign GEN_49 = reg_tselect ? reg_bp_1_control_tmatch : reg_bp_0_control_tmatch;
  assign GEN_50 = reg_tselect ? reg_bp_1_control_m : reg_bp_0_control_m;
  assign GEN_51 = reg_tselect ? reg_bp_1_control_h : reg_bp_0_control_h;
  assign GEN_52 = reg_tselect ? reg_bp_1_control_s : reg_bp_0_control_s;
  assign GEN_53 = reg_tselect ? reg_bp_1_control_u : reg_bp_0_control_u;
  assign GEN_54 = reg_tselect ? reg_bp_1_control_x : reg_bp_0_control_x;
  assign GEN_55 = reg_tselect ? reg_bp_1_control_w : reg_bp_0_control_w;
  assign GEN_56 = reg_tselect ? reg_bp_1_control_r : reg_bp_0_control_r;
  assign GEN_57 = reg_tselect ? reg_bp_1_address : reg_bp_0_address;
  assign GEN_1_control_ttype = GEN_42;
  assign GEN_1_control_dmode = GEN_43;
  assign GEN_1_control_maskmax = GEN_44;
  assign GEN_1_control_reserved = GEN_45;
  assign GEN_1_control_action = GEN_46;
  assign GEN_1_control_chain = GEN_47;
  assign GEN_1_control_zero = GEN_48;
  assign GEN_1_control_tmatch = GEN_49;
  assign GEN_1_control_m = GEN_50;
  assign GEN_1_control_h = GEN_51;
  assign GEN_1_control_s = GEN_52;
  assign GEN_1_control_u = GEN_53;
  assign GEN_1_control_x = GEN_54;
  assign GEN_1_control_w = GEN_55;
  assign GEN_1_control_r = GEN_56;
  assign GEN_1_address = GEN_57;
  assign T_5885 = {GEN_0_control_x,GEN_1_control_w};
  assign GEN_2_control_ttype = GEN_42;
  assign GEN_2_control_dmode = GEN_43;
  assign GEN_2_control_maskmax = GEN_44;
  assign GEN_2_control_reserved = GEN_45;
  assign GEN_2_control_action = GEN_46;
  assign GEN_2_control_chain = GEN_47;
  assign GEN_2_control_zero = GEN_48;
  assign GEN_2_control_tmatch = GEN_49;
  assign GEN_2_control_m = GEN_50;
  assign GEN_2_control_h = GEN_51;
  assign GEN_2_control_s = GEN_52;
  assign GEN_2_control_u = GEN_53;
  assign GEN_2_control_x = GEN_54;
  assign GEN_2_control_w = GEN_55;
  assign GEN_2_control_r = GEN_56;
  assign GEN_2_address = GEN_57;
  assign T_5886 = {T_5885,GEN_2_control_r};
  assign GEN_3_control_ttype = GEN_42;
  assign GEN_3_control_dmode = GEN_43;
  assign GEN_3_control_maskmax = GEN_44;
  assign GEN_3_control_reserved = GEN_45;
  assign GEN_3_control_action = GEN_46;
  assign GEN_3_control_chain = GEN_47;
  assign GEN_3_control_zero = GEN_48;
  assign GEN_3_control_tmatch = GEN_49;
  assign GEN_3_control_m = GEN_50;
  assign GEN_3_control_h = GEN_51;
  assign GEN_3_control_s = GEN_52;
  assign GEN_3_control_u = GEN_53;
  assign GEN_3_control_x = GEN_54;
  assign GEN_3_control_w = GEN_55;
  assign GEN_3_control_r = GEN_56;
  assign GEN_3_address = GEN_57;
  assign GEN_4_control_ttype = GEN_42;
  assign GEN_4_control_dmode = GEN_43;
  assign GEN_4_control_maskmax = GEN_44;
  assign GEN_4_control_reserved = GEN_45;
  assign GEN_4_control_action = GEN_46;
  assign GEN_4_control_chain = GEN_47;
  assign GEN_4_control_zero = GEN_48;
  assign GEN_4_control_tmatch = GEN_49;
  assign GEN_4_control_m = GEN_50;
  assign GEN_4_control_h = GEN_51;
  assign GEN_4_control_s = GEN_52;
  assign GEN_4_control_u = GEN_53;
  assign GEN_4_control_x = GEN_54;
  assign GEN_4_control_w = GEN_55;
  assign GEN_4_control_r = GEN_56;
  assign GEN_4_address = GEN_57;
  assign T_5887 = {GEN_3_control_s,GEN_4_control_u};
  assign GEN_5_control_ttype = GEN_42;
  assign GEN_5_control_dmode = GEN_43;
  assign GEN_5_control_maskmax = GEN_44;
  assign GEN_5_control_reserved = GEN_45;
  assign GEN_5_control_action = GEN_46;
  assign GEN_5_control_chain = GEN_47;
  assign GEN_5_control_zero = GEN_48;
  assign GEN_5_control_tmatch = GEN_49;
  assign GEN_5_control_m = GEN_50;
  assign GEN_5_control_h = GEN_51;
  assign GEN_5_control_s = GEN_52;
  assign GEN_5_control_u = GEN_53;
  assign GEN_5_control_x = GEN_54;
  assign GEN_5_control_w = GEN_55;
  assign GEN_5_control_r = GEN_56;
  assign GEN_5_address = GEN_57;
  assign GEN_6_control_ttype = GEN_42;
  assign GEN_6_control_dmode = GEN_43;
  assign GEN_6_control_maskmax = GEN_44;
  assign GEN_6_control_reserved = GEN_45;
  assign GEN_6_control_action = GEN_46;
  assign GEN_6_control_chain = GEN_47;
  assign GEN_6_control_zero = GEN_48;
  assign GEN_6_control_tmatch = GEN_49;
  assign GEN_6_control_m = GEN_50;
  assign GEN_6_control_h = GEN_51;
  assign GEN_6_control_s = GEN_52;
  assign GEN_6_control_u = GEN_53;
  assign GEN_6_control_x = GEN_54;
  assign GEN_6_control_w = GEN_55;
  assign GEN_6_control_r = GEN_56;
  assign GEN_6_address = GEN_57;
  assign T_5888 = {GEN_5_control_m,GEN_6_control_h};
  assign T_5889 = {T_5888,T_5887};
  assign T_5890 = {T_5889,T_5886};
  assign GEN_7_control_ttype = GEN_42;
  assign GEN_7_control_dmode = GEN_43;
  assign GEN_7_control_maskmax = GEN_44;
  assign GEN_7_control_reserved = GEN_45;
  assign GEN_7_control_action = GEN_46;
  assign GEN_7_control_chain = GEN_47;
  assign GEN_7_control_zero = GEN_48;
  assign GEN_7_control_tmatch = GEN_49;
  assign GEN_7_control_m = GEN_50;
  assign GEN_7_control_h = GEN_51;
  assign GEN_7_control_s = GEN_52;
  assign GEN_7_control_u = GEN_53;
  assign GEN_7_control_x = GEN_54;
  assign GEN_7_control_w = GEN_55;
  assign GEN_7_control_r = GEN_56;
  assign GEN_7_address = GEN_57;
  assign GEN_8_control_ttype = GEN_42;
  assign GEN_8_control_dmode = GEN_43;
  assign GEN_8_control_maskmax = GEN_44;
  assign GEN_8_control_reserved = GEN_45;
  assign GEN_8_control_action = GEN_46;
  assign GEN_8_control_chain = GEN_47;
  assign GEN_8_control_zero = GEN_48;
  assign GEN_8_control_tmatch = GEN_49;
  assign GEN_8_control_m = GEN_50;
  assign GEN_8_control_h = GEN_51;
  assign GEN_8_control_s = GEN_52;
  assign GEN_8_control_u = GEN_53;
  assign GEN_8_control_x = GEN_54;
  assign GEN_8_control_w = GEN_55;
  assign GEN_8_control_r = GEN_56;
  assign GEN_8_address = GEN_57;
  assign T_5891 = {GEN_7_control_zero,GEN_8_control_tmatch};
  assign GEN_9_control_ttype = GEN_42;
  assign GEN_9_control_dmode = GEN_43;
  assign GEN_9_control_maskmax = GEN_44;
  assign GEN_9_control_reserved = GEN_45;
  assign GEN_9_control_action = GEN_46;
  assign GEN_9_control_chain = GEN_47;
  assign GEN_9_control_zero = GEN_48;
  assign GEN_9_control_tmatch = GEN_49;
  assign GEN_9_control_m = GEN_50;
  assign GEN_9_control_h = GEN_51;
  assign GEN_9_control_s = GEN_52;
  assign GEN_9_control_u = GEN_53;
  assign GEN_9_control_x = GEN_54;
  assign GEN_9_control_w = GEN_55;
  assign GEN_9_control_r = GEN_56;
  assign GEN_9_address = GEN_57;
  assign GEN_10_control_ttype = GEN_42;
  assign GEN_10_control_dmode = GEN_43;
  assign GEN_10_control_maskmax = GEN_44;
  assign GEN_10_control_reserved = GEN_45;
  assign GEN_10_control_action = GEN_46;
  assign GEN_10_control_chain = GEN_47;
  assign GEN_10_control_zero = GEN_48;
  assign GEN_10_control_tmatch = GEN_49;
  assign GEN_10_control_m = GEN_50;
  assign GEN_10_control_h = GEN_51;
  assign GEN_10_control_s = GEN_52;
  assign GEN_10_control_u = GEN_53;
  assign GEN_10_control_x = GEN_54;
  assign GEN_10_control_w = GEN_55;
  assign GEN_10_control_r = GEN_56;
  assign GEN_10_address = GEN_57;
  assign T_5892 = {GEN_9_control_action,GEN_10_control_chain};
  assign T_5893 = {T_5892,T_5891};
  assign GEN_11_control_ttype = GEN_42;
  assign GEN_11_control_dmode = GEN_43;
  assign GEN_11_control_maskmax = GEN_44;
  assign GEN_11_control_reserved = GEN_45;
  assign GEN_11_control_action = GEN_46;
  assign GEN_11_control_chain = GEN_47;
  assign GEN_11_control_zero = GEN_48;
  assign GEN_11_control_tmatch = GEN_49;
  assign GEN_11_control_m = GEN_50;
  assign GEN_11_control_h = GEN_51;
  assign GEN_11_control_s = GEN_52;
  assign GEN_11_control_u = GEN_53;
  assign GEN_11_control_x = GEN_54;
  assign GEN_11_control_w = GEN_55;
  assign GEN_11_control_r = GEN_56;
  assign GEN_11_address = GEN_57;
  assign GEN_12_control_ttype = GEN_42;
  assign GEN_12_control_dmode = GEN_43;
  assign GEN_12_control_maskmax = GEN_44;
  assign GEN_12_control_reserved = GEN_45;
  assign GEN_12_control_action = GEN_46;
  assign GEN_12_control_chain = GEN_47;
  assign GEN_12_control_zero = GEN_48;
  assign GEN_12_control_tmatch = GEN_49;
  assign GEN_12_control_m = GEN_50;
  assign GEN_12_control_h = GEN_51;
  assign GEN_12_control_s = GEN_52;
  assign GEN_12_control_u = GEN_53;
  assign GEN_12_control_x = GEN_54;
  assign GEN_12_control_w = GEN_55;
  assign GEN_12_control_r = GEN_56;
  assign GEN_12_address = GEN_57;
  assign T_5894 = {GEN_11_control_maskmax,GEN_12_control_reserved};
  assign GEN_13_control_ttype = GEN_42;
  assign GEN_13_control_dmode = GEN_43;
  assign GEN_13_control_maskmax = GEN_44;
  assign GEN_13_control_reserved = GEN_45;
  assign GEN_13_control_action = GEN_46;
  assign GEN_13_control_chain = GEN_47;
  assign GEN_13_control_zero = GEN_48;
  assign GEN_13_control_tmatch = GEN_49;
  assign GEN_13_control_m = GEN_50;
  assign GEN_13_control_h = GEN_51;
  assign GEN_13_control_s = GEN_52;
  assign GEN_13_control_u = GEN_53;
  assign GEN_13_control_x = GEN_54;
  assign GEN_13_control_w = GEN_55;
  assign GEN_13_control_r = GEN_56;
  assign GEN_13_address = GEN_57;
  assign GEN_14_control_ttype = GEN_42;
  assign GEN_14_control_dmode = GEN_43;
  assign GEN_14_control_maskmax = GEN_44;
  assign GEN_14_control_reserved = GEN_45;
  assign GEN_14_control_action = GEN_46;
  assign GEN_14_control_chain = GEN_47;
  assign GEN_14_control_zero = GEN_48;
  assign GEN_14_control_tmatch = GEN_49;
  assign GEN_14_control_m = GEN_50;
  assign GEN_14_control_h = GEN_51;
  assign GEN_14_control_s = GEN_52;
  assign GEN_14_control_u = GEN_53;
  assign GEN_14_control_x = GEN_54;
  assign GEN_14_control_w = GEN_55;
  assign GEN_14_control_r = GEN_56;
  assign GEN_14_address = GEN_57;
  assign T_5895 = {GEN_13_control_ttype,GEN_14_control_dmode};
  assign T_5896 = {T_5895,T_5894};
  assign T_5897 = {T_5896,T_5893};
  assign T_5898 = {T_5897,T_5890};
  assign GEN_15_control_ttype = GEN_42;
  assign GEN_15_control_dmode = GEN_43;
  assign GEN_15_control_maskmax = GEN_44;
  assign GEN_15_control_reserved = GEN_45;
  assign GEN_15_control_action = GEN_46;
  assign GEN_15_control_chain = GEN_47;
  assign GEN_15_control_zero = GEN_48;
  assign GEN_15_control_tmatch = GEN_49;
  assign GEN_15_control_m = GEN_50;
  assign GEN_15_control_h = GEN_51;
  assign GEN_15_control_s = GEN_52;
  assign GEN_15_control_u = GEN_53;
  assign GEN_15_control_x = GEN_54;
  assign GEN_15_control_w = GEN_55;
  assign GEN_15_control_r = GEN_56;
  assign GEN_15_address = GEN_57;
  assign T_5916 = GEN_15_address[38];
  assign T_5920 = T_5916 ? 25'h1ffffff : 25'h0;
  assign GEN_16_control_ttype = GEN_42;
  assign GEN_16_control_dmode = GEN_43;
  assign GEN_16_control_maskmax = GEN_44;
  assign GEN_16_control_reserved = GEN_45;
  assign GEN_16_control_action = GEN_46;
  assign GEN_16_control_chain = GEN_47;
  assign GEN_16_control_zero = GEN_48;
  assign GEN_16_control_tmatch = GEN_49;
  assign GEN_16_control_m = GEN_50;
  assign GEN_16_control_h = GEN_51;
  assign GEN_16_control_s = GEN_52;
  assign GEN_16_control_u = GEN_53;
  assign GEN_16_control_x = GEN_54;
  assign GEN_16_control_w = GEN_55;
  assign GEN_16_control_r = GEN_56;
  assign GEN_16_address = GEN_57;
  assign T_5921 = {T_5920,GEN_16_address};
  assign T_5926 = reg_mepc[39];
  assign T_5930 = T_5926 ? 24'hffffff : 24'h0;
  assign T_5931 = {T_5930,reg_mepc};
  assign T_5932 = reg_mbadaddr[39];
  assign T_5936 = T_5932 ? 24'hffffff : 24'h0;
  assign T_5937 = {T_5936,reg_mbadaddr};
  assign T_5938 = {reg_dcsr_step,reg_dcsr_prv};
  assign T_5939 = {reg_dcsr_zero1,reg_dcsr_halt};
  assign T_5940 = {T_5939,T_5938};
  assign T_5941 = {reg_dcsr_cause,reg_dcsr_debugint};
  assign T_5942 = {reg_dcsr_stopcycle,reg_dcsr_stoptime};
  assign T_5943 = {T_5942,T_5941};
  assign T_5944 = {T_5943,T_5940};
  assign T_5945 = {reg_dcsr_ebreaku,reg_dcsr_zero2};
  assign T_5946 = {reg_dcsr_ebreakh,reg_dcsr_ebreaks};
  assign T_5947 = {T_5946,T_5945};
  assign T_5948 = {reg_dcsr_zero3,reg_dcsr_ebreakm};
  assign T_5949 = {reg_dcsr_xdebugver,reg_dcsr_ndreset};
  assign T_5950 = {T_5949,reg_dcsr_fullreset};
  assign T_5951 = {T_5950,T_5948};
  assign T_5952 = {T_5951,T_5947};
  assign T_5953 = {T_5952,T_5944};
  assign T_5958 = io_rw_addr == 12'h7a0;
  assign T_5960 = io_rw_addr == 12'h7a1;
  assign T_5962 = io_rw_addr == 12'h7a2;
  assign T_5964 = io_rw_addr == 12'hf13;
  assign T_5966 = io_rw_addr == 12'hf12;
  assign T_5968 = io_rw_addr == 12'hf11;
  assign T_5970 = io_rw_addr == 12'hb00;
  assign T_5972 = io_rw_addr == 12'hb02;
  assign T_5974 = io_rw_addr == 12'h301;
  assign T_5976 = io_rw_addr == 12'h300;
  assign T_5978 = io_rw_addr == 12'h305;
  assign T_5980 = io_rw_addr == 12'h344;
  assign T_5982 = io_rw_addr == 12'h304;
  assign T_5984 = io_rw_addr == 12'h303;
  assign T_5986 = io_rw_addr == 12'h302;
  assign T_5988 = io_rw_addr == 12'h340;
  assign T_5990 = io_rw_addr == 12'h341;
  assign T_5992 = io_rw_addr == 12'h343;
  assign T_5994 = io_rw_addr == 12'h342;
  assign T_5996 = io_rw_addr == 12'hf14;
  assign T_5998 = io_rw_addr == 12'h7b0;
  assign T_6000 = io_rw_addr == 12'h7b1;
  assign T_6002 = io_rw_addr == 12'h7b2;
  assign T_6004 = io_rw_addr == 12'h323;
  assign T_6006 = io_rw_addr == 12'hb03;
  assign T_6008 = io_rw_addr == 12'h324;
  assign T_6010 = io_rw_addr == 12'hb04;
  assign T_6012 = io_rw_addr == 12'h325;
  assign T_6014 = io_rw_addr == 12'hb05;
  assign T_6016 = io_rw_addr == 12'h326;
  assign T_6018 = io_rw_addr == 12'hb06;
  assign T_6020 = io_rw_addr == 12'h327;
  assign T_6022 = io_rw_addr == 12'hb07;
  assign T_6024 = io_rw_addr == 12'h328;
  assign T_6026 = io_rw_addr == 12'hb08;
  assign T_6028 = io_rw_addr == 12'h329;
  assign T_6030 = io_rw_addr == 12'hb09;
  assign T_6032 = io_rw_addr == 12'h32a;
  assign T_6034 = io_rw_addr == 12'hb0a;
  assign T_6036 = io_rw_addr == 12'h32b;
  assign T_6038 = io_rw_addr == 12'hb0b;
  assign T_6040 = io_rw_addr == 12'h32c;
  assign T_6042 = io_rw_addr == 12'hb0c;
  assign T_6044 = io_rw_addr == 12'h32d;
  assign T_6046 = io_rw_addr == 12'hb0d;
  assign T_6048 = io_rw_addr == 12'h32e;
  assign T_6050 = io_rw_addr == 12'hb0e;
  assign T_6052 = io_rw_addr == 12'h32f;
  assign T_6054 = io_rw_addr == 12'hb0f;
  assign T_6056 = io_rw_addr == 12'h330;
  assign T_6058 = io_rw_addr == 12'hb10;
  assign T_6060 = io_rw_addr == 12'h331;
  assign T_6062 = io_rw_addr == 12'hb11;
  assign T_6064 = io_rw_addr == 12'h332;
  assign T_6066 = io_rw_addr == 12'hb12;
  assign T_6068 = io_rw_addr == 12'h333;
  assign T_6070 = io_rw_addr == 12'hb13;
  assign T_6072 = io_rw_addr == 12'h334;
  assign T_6074 = io_rw_addr == 12'hb14;
  assign T_6076 = io_rw_addr == 12'h335;
  assign T_6078 = io_rw_addr == 12'hb15;
  assign T_6080 = io_rw_addr == 12'h336;
  assign T_6082 = io_rw_addr == 12'hb16;
  assign T_6084 = io_rw_addr == 12'h337;
  assign T_6086 = io_rw_addr == 12'hb17;
  assign T_6088 = io_rw_addr == 12'h338;
  assign T_6090 = io_rw_addr == 12'hb18;
  assign T_6092 = io_rw_addr == 12'h339;
  assign T_6094 = io_rw_addr == 12'hb19;
  assign T_6096 = io_rw_addr == 12'h33a;
  assign T_6098 = io_rw_addr == 12'hb1a;
  assign T_6100 = io_rw_addr == 12'h33b;
  assign T_6102 = io_rw_addr == 12'hb1b;
  assign T_6104 = io_rw_addr == 12'h33c;
  assign T_6106 = io_rw_addr == 12'hb1c;
  assign T_6108 = io_rw_addr == 12'h33d;
  assign T_6110 = io_rw_addr == 12'hb1d;
  assign T_6112 = io_rw_addr == 12'h33e;
  assign T_6114 = io_rw_addr == 12'hb1e;
  assign T_6116 = io_rw_addr == 12'h33f;
  assign T_6118 = io_rw_addr == 12'hb1f;
  assign T_6119 = T_5958 | T_5960;
  assign T_6120 = T_6119 | T_5962;
  assign T_6121 = T_6120 | T_5964;
  assign T_6122 = T_6121 | T_5966;
  assign T_6123 = T_6122 | T_5968;
  assign T_6124 = T_6123 | T_5970;
  assign T_6125 = T_6124 | T_5972;
  assign T_6126 = T_6125 | T_5974;
  assign T_6127 = T_6126 | T_5976;
  assign T_6128 = T_6127 | T_5978;
  assign T_6129 = T_6128 | T_5980;
  assign T_6130 = T_6129 | T_5982;
  assign T_6131 = T_6130 | T_5984;
  assign T_6132 = T_6131 | T_5986;
  assign T_6133 = T_6132 | T_5988;
  assign T_6134 = T_6133 | T_5990;
  assign T_6135 = T_6134 | T_5992;
  assign T_6136 = T_6135 | T_5994;
  assign T_6137 = T_6136 | T_5996;
  assign T_6138 = T_6137 | T_5998;
  assign T_6139 = T_6138 | T_6000;
  assign T_6140 = T_6139 | T_6002;
  assign T_6141 = T_6140 | T_6004;
  assign T_6142 = T_6141 | T_6006;
  assign T_6143 = T_6142 | T_6008;
  assign T_6144 = T_6143 | T_6010;
  assign T_6145 = T_6144 | T_6012;
  assign T_6146 = T_6145 | T_6014;
  assign T_6147 = T_6146 | T_6016;
  assign T_6148 = T_6147 | T_6018;
  assign T_6149 = T_6148 | T_6020;
  assign T_6150 = T_6149 | T_6022;
  assign T_6151 = T_6150 | T_6024;
  assign T_6152 = T_6151 | T_6026;
  assign T_6153 = T_6152 | T_6028;
  assign T_6154 = T_6153 | T_6030;
  assign T_6155 = T_6154 | T_6032;
  assign T_6156 = T_6155 | T_6034;
  assign T_6157 = T_6156 | T_6036;
  assign T_6158 = T_6157 | T_6038;
  assign T_6159 = T_6158 | T_6040;
  assign T_6160 = T_6159 | T_6042;
  assign T_6161 = T_6160 | T_6044;
  assign T_6162 = T_6161 | T_6046;
  assign T_6163 = T_6162 | T_6048;
  assign T_6164 = T_6163 | T_6050;
  assign T_6165 = T_6164 | T_6052;
  assign T_6166 = T_6165 | T_6054;
  assign T_6167 = T_6166 | T_6056;
  assign T_6168 = T_6167 | T_6058;
  assign T_6169 = T_6168 | T_6060;
  assign T_6170 = T_6169 | T_6062;
  assign T_6171 = T_6170 | T_6064;
  assign T_6172 = T_6171 | T_6066;
  assign T_6173 = T_6172 | T_6068;
  assign T_6174 = T_6173 | T_6070;
  assign T_6175 = T_6174 | T_6072;
  assign T_6176 = T_6175 | T_6074;
  assign T_6177 = T_6176 | T_6076;
  assign T_6178 = T_6177 | T_6078;
  assign T_6179 = T_6178 | T_6080;
  assign T_6180 = T_6179 | T_6082;
  assign T_6181 = T_6180 | T_6084;
  assign T_6182 = T_6181 | T_6086;
  assign T_6183 = T_6182 | T_6088;
  assign T_6184 = T_6183 | T_6090;
  assign T_6185 = T_6184 | T_6092;
  assign T_6186 = T_6185 | T_6094;
  assign T_6187 = T_6186 | T_6096;
  assign T_6188 = T_6187 | T_6098;
  assign T_6189 = T_6188 | T_6100;
  assign T_6190 = T_6189 | T_6102;
  assign T_6191 = T_6190 | T_6104;
  assign T_6192 = T_6191 | T_6106;
  assign T_6193 = T_6192 | T_6108;
  assign T_6194 = T_6193 | T_6110;
  assign T_6195 = T_6194 | T_6112;
  assign T_6196 = T_6195 | T_6114;
  assign T_6197 = T_6196 | T_6116;
  assign addr_valid = T_6197 | T_6118;
  assign csr_addr_priv = io_rw_addr[9:8];
  assign T_6216 = io_rw_addr & 12'h90;
  assign T_6218 = T_6216 == 12'h90;
  assign T_6220 = T_6218 == 1'h0;
  assign T_6221 = reg_mstatus_prv >= csr_addr_priv;
  assign T_6222 = T_6220 & T_6221;
  assign priv_sufficient = reg_debug | T_6222;
  assign T_6223 = io_rw_addr[11:10];
  assign T_6224 = ~ T_6223;
  assign read_only = T_6224 == 2'h0;
  assign T_6226 = cpu_wen & priv_sufficient;
  assign T_6228 = read_only == 1'h0;
  assign wen = T_6226 & T_6228;
  assign T_6229 = io_rw_cmd == 3'h2;
  assign T_6230 = io_rw_cmd == 3'h3;
  assign T_6231 = T_6229 | T_6230;
  assign T_6233 = T_6231 ? io_rw_rdata : 64'h0;
  assign T_6234 = io_rw_cmd != 3'h3;
  assign T_6236 = T_6234 ? io_rw_wdata : 64'h0;
  assign T_6237 = T_6233 | T_6236;
  assign T_6240 = T_6230 ? io_rw_wdata : 64'h0;
  assign T_6241 = ~ T_6240;
  assign wdata = T_6237 & T_6241;
  assign do_system_insn = priv_sufficient & system_insn;
  assign T_6243 = io_rw_addr[2:0];
  assign opcode = 8'h1 << T_6243;
  assign T_6244 = opcode[0];
  assign insn_call = do_system_insn & T_6244;
  assign T_6245 = opcode[1];
  assign insn_break = do_system_insn & T_6245;
  assign T_6246 = opcode[2];
  assign insn_ret = do_system_insn & T_6246;
  assign T_6247 = opcode[4];
  assign insn_sfence_vm = do_system_insn & T_6247;
  assign T_6248 = opcode[5];
  assign insn_wfi = do_system_insn & T_6248;
  assign T_6249 = cpu_wen & read_only;
  assign T_6251 = priv_sufficient == 1'h0;
  assign T_6253 = addr_valid == 1'h0;
  assign T_6254 = T_6251 | T_6253;
  assign T_6265 = cpu_ren & T_6254;
  assign T_6266 = T_6249 | T_6265;
  assign T_6269 = system_insn & T_6251;
  assign T_6270 = T_6266 | T_6269;
  assign T_6271 = T_6270 | insn_call;
  assign T_6272 = T_6271 | insn_break;
  assign GEN_314 = insn_wfi ? 1'h1 : reg_wfi;
  assign T_6275 = pending_interrupts != 64'h0;
  assign GEN_315 = T_6275 ? 1'h0 : GEN_314;
  assign T_6278 = io_csr_xcpt == 1'h0;
  assign GEN_3 = {{2'd0}, reg_mstatus_prv};
  assign T_6280 = GEN_3 + 4'h8;
  assign T_6281 = T_6280[3:0];
  assign T_6284 = insn_break ? 2'h3 : 2'h2;
  assign T_6285 = insn_call ? T_6281 : {{2'd0}, T_6284};
  assign cause = T_6278 ? io_cause : {{60'd0}, T_6285};
  assign cause_lsbs = cause[5:0];
  assign T_6286 = cause[63];
  assign T_6288 = cause_lsbs == 6'hd;
  assign causeIsDebugInt = T_6286 & T_6288;
  assign T_6291 = T_6286 == 1'h0;
  assign causeIsDebugTrigger = T_6291 & T_6288;
  assign T_6297 = T_6291 & insn_break;
  assign T_6298 = {reg_dcsr_ebreaks,reg_dcsr_ebreaku};
  assign T_6299 = {reg_dcsr_ebreakm,reg_dcsr_ebreakh};
  assign T_6300 = {T_6299,T_6298};
  assign T_6301 = T_6300 >> reg_mstatus_prv;
  assign T_6302 = T_6301[0];
  assign causeIsDebugBreak = T_6297 & T_6302;
  assign T_6304 = reg_singleStepped | causeIsDebugInt;
  assign T_6305 = T_6304 | causeIsDebugTrigger;
  assign T_6306 = T_6305 | causeIsDebugBreak;
  assign T_6307 = T_6306 | reg_debug;
  assign debugTVec = reg_debug ? 12'h808 : 12'h800;
  assign T_6322 = {{8'd0}, reg_mtvec};
  assign tvec = T_6307 ? {{28'd0}, debugTVec} : T_6322;
  assign epc = T_6218 ? reg_dpc : reg_mepc;
  assign T_6329 = exception ? tvec : epc;
  assign T_6332 = reg_dcsr_step & T_5613;
  assign T_6333 = ~ io_status_fs;
  assign T_6335 = T_6333 == 2'h0;
  assign T_6336 = ~ io_status_xs;
  assign T_6338 = T_6336 == 2'h0;
  assign T_6339 = T_6335 | T_6338;
  assign T_6340 = ~ io_pc;
  assign T_6342 = T_6340 | 40'h1;
  assign T_6343 = ~ T_6342;
  assign T_6344 = read_mstatus >> reg_mstatus_prv;
  assign T_6345 = T_6344[0];
  assign T_6353 = cause == 64'h3;
  assign T_6354 = cause == 64'h4;
  assign T_6355 = cause == 64'h6;
  assign T_6356 = cause == 64'h0;
  assign T_6357 = cause == 64'h5;
  assign T_6358 = cause == 64'h7;
  assign T_6359 = cause == 64'h1;
  assign T_6360 = T_6353 | T_6354;
  assign T_6361 = T_6360 | T_6355;
  assign T_6362 = T_6361 | T_6356;
  assign T_6363 = T_6362 | T_6357;
  assign T_6364 = T_6363 | T_6358;
  assign T_6365 = T_6364 | T_6359;
  assign T_6371 = causeIsDebugTrigger ? 2'h2 : 2'h1;
  assign T_6372 = causeIsDebugInt ? 2'h3 : T_6371;
  assign T_6373 = reg_singleStepped ? 3'h4 : {{1'd0}, T_6372};
  assign GEN_316 = T_6307 ? 1'h1 : reg_debug;
  assign GEN_317 = T_6307 ? T_6343 : reg_dpc;
  assign GEN_318 = T_6307 ? T_6373 : reg_dcsr_cause;
  assign GEN_319 = T_6307 ? 2'h3 : reg_dcsr_prv;
  assign T_6376 = T_6307 == 1'h0;
  assign GEN_325 = {{1'd0}, reg_mstatus_spp};
  assign GEN_328 = T_6365 ? io_badaddr : reg_mbadaddr;
  assign GEN_329 = T_6376 ? T_6343 : reg_mepc;
  assign GEN_330 = T_6376 ? cause : reg_mcause;
  assign GEN_331 = T_6376 ? GEN_328 : reg_mbadaddr;
  assign GEN_332 = T_6376 ? T_6345 : reg_mstatus_mpie;
  assign GEN_333 = T_6376 ? 2'h3 : reg_mstatus_mpp;
  assign GEN_334 = T_6376 ? 1'h0 : reg_mstatus_mie;
  assign GEN_335 = T_6376 ? 2'h3 : reg_mstatus_prv;
  assign GEN_336 = exception ? GEN_316 : reg_debug;
  assign GEN_337 = exception ? GEN_317 : reg_dpc;
  assign GEN_338 = exception ? GEN_318 : reg_dcsr_cause;
  assign GEN_339 = exception ? GEN_319 : reg_dcsr_prv;
  assign GEN_344 = exception ? GEN_325 : {{1'd0}, reg_mstatus_spp};
  assign GEN_346 = exception ? GEN_335 : reg_mstatus_prv;
  assign GEN_347 = exception ? GEN_329 : reg_mepc;
  assign GEN_348 = exception ? GEN_330 : reg_mcause;
  assign GEN_349 = exception ? GEN_331 : reg_mbadaddr;
  assign GEN_350 = exception ? GEN_332 : reg_mstatus_mpie;
  assign GEN_351 = exception ? GEN_333 : reg_mstatus_mpp;
  assign GEN_352 = exception ? GEN_334 : reg_mstatus_mie;
  assign GEN_358 = T_6218 ? reg_dcsr_prv : GEN_346;
  assign GEN_359 = T_6218 ? 1'h0 : GEN_336;
  assign T_6405 = reg_mstatus_mpp[1];
  assign GEN_360 = T_6405 ? reg_mstatus_mpie : GEN_352;
  assign GEN_362 = T_6220 ? GEN_360 : GEN_352;
  assign GEN_364 = T_6220 ? 1'h0 : GEN_350;
  assign GEN_365 = T_6220 ? 2'h3 : GEN_351;
  assign GEN_366 = T_6220 ? reg_mstatus_mpp : GEN_358;
  assign GEN_370 = insn_ret ? GEN_366 : GEN_346;
  assign GEN_371 = insn_ret ? GEN_359 : GEN_336;
  assign GEN_372 = insn_ret ? GEN_362 : GEN_352;
  assign GEN_373 = insn_ret ? GEN_364 : GEN_350;
  assign GEN_374 = insn_ret ? GEN_365 : GEN_351;
  assign T_6415 = io_exception + io_csr_xcpt;
  assign GEN_4 = {{1'd0}, insn_ret};
  assign T_6416 = GEN_4 + T_6415;
  assign T_6418 = T_6416 <= 3'h1;
  assign T_6419 = T_6418 | reset;
  assign T_6421 = T_6419 == 1'h0;
  assign T_6423 = T_5958 ? reg_tselect : 1'h0;
  assign T_6425 = T_5960 ? T_5898 : 64'h0;
  assign T_6427 = T_5962 ? T_5921 : 64'h0;
  assign T_6435 = T_5970 ? T_5586 : 64'h0;
  assign T_6437 = T_5972 ? T_5575 : 64'h0;
  assign T_6439 = T_5974 ? 64'h8000000000001101 : 64'h0;
  assign T_6441 = T_5976 ? read_mstatus : 64'h0;
  assign T_6443 = T_5978 ? reg_mtvec : 32'h0;
  assign T_6445 = T_5980 ? read_mip : 13'h0;
  assign T_6447 = T_5982 ? reg_mie : 64'h0;
  assign T_6449 = T_5984 ? reg_mideleg : 64'h0;
  assign T_6451 = T_5986 ? reg_medeleg : 64'h0;
  assign T_6453 = T_5988 ? reg_mscratch : 64'h0;
  assign T_6455 = T_5990 ? T_5931 : 64'h0;
  assign T_6457 = T_5992 ? T_5937 : 64'h0;
  assign T_6459 = T_5994 ? reg_mcause : 64'h0;
  assign T_6461 = T_5996 ? io_prci_id : 1'h0;
  assign T_6463 = T_5998 ? T_5953 : 32'h0;
  assign T_6465 = T_6000 ? reg_dpc : 40'h0;
  assign T_6467 = T_6002 ? reg_dscratch : 64'h0;
  assign GEN_5 = {{63'd0}, T_6423};
  assign T_6585 = GEN_5 | T_6425;
  assign T_6586 = T_6585 | T_6427;
  assign T_6590 = T_6586 | T_6435;
  assign T_6591 = T_6590 | T_6437;
  assign T_6592 = T_6591 | T_6439;
  assign T_6593 = T_6592 | T_6441;
  assign GEN_6 = {{32'd0}, T_6443};
  assign T_6594 = T_6593 | GEN_6;
  assign GEN_7 = {{51'd0}, T_6445};
  assign T_6595 = T_6594 | GEN_7;
  assign T_6596 = T_6595 | T_6447;
  assign T_6597 = T_6596 | T_6449;
  assign T_6598 = T_6597 | T_6451;
  assign T_6599 = T_6598 | T_6453;
  assign T_6600 = T_6599 | T_6455;
  assign T_6601 = T_6600 | T_6457;
  assign T_6602 = T_6601 | T_6459;
  assign GEN_8 = {{63'd0}, T_6461};
  assign T_6603 = T_6602 | GEN_8;
  assign GEN_9 = {{32'd0}, T_6463};
  assign T_6604 = T_6603 | GEN_9;
  assign GEN_10 = {{24'd0}, T_6465};
  assign T_6605 = T_6604 | GEN_10;
  assign T_6606 = T_6605 | T_6467;
  assign T_6665 = T_6606;
  assign T_6666 = reg_fflags | io_fcsr_flags_bits;
  assign GEN_375 = io_fcsr_flags_valid ? T_6666 : reg_fflags;
  assign T_6717_debug = T_6767;
  assign T_6717_prv = T_6766;
  assign T_6717_sd = T_6765;
  assign T_6717_zero3 = T_6764;
  assign T_6717_sd_rv32 = T_6763;
  assign T_6717_zero2 = T_6762;
  assign T_6717_vm = T_6761;
  assign T_6717_zero1 = T_6760;
  assign T_6717_mxr = T_6759;
  assign T_6717_pum = T_6758;
  assign T_6717_mprv = T_6757;
  assign T_6717_xs = T_6756;
  assign T_6717_fs = T_6755;
  assign T_6717_mpp = T_6754;
  assign T_6717_hpp = T_6753;
  assign T_6717_spp = T_6752;
  assign T_6717_mpie = T_6751;
  assign T_6717_hpie = T_6750;
  assign T_6717_spie = T_6749;
  assign T_6717_upie = T_6748;
  assign T_6717_mie = T_6747;
  assign T_6717_hie = T_6746;
  assign T_6717_sie = T_6745;
  assign T_6717_uie = T_6744;
  assign T_6743 = {{3'd0}, wdata};
  assign T_6744 = T_6743[0];
  assign T_6745 = T_6743[1];
  assign T_6746 = T_6743[2];
  assign T_6747 = T_6743[3];
  assign T_6748 = T_6743[4];
  assign T_6749 = T_6743[5];
  assign T_6750 = T_6743[6];
  assign T_6751 = T_6743[7];
  assign T_6752 = T_6743[8];
  assign T_6753 = T_6743[10:9];
  assign T_6754 = T_6743[12:11];
  assign T_6755 = T_6743[14:13];
  assign T_6756 = T_6743[16:15];
  assign T_6757 = T_6743[17];
  assign T_6758 = T_6743[18];
  assign T_6759 = T_6743[19];
  assign T_6760 = T_6743[23:20];
  assign T_6761 = T_6743[28:24];
  assign T_6762 = T_6743[30:29];
  assign T_6763 = T_6743[31];
  assign T_6764 = T_6743[62:32];
  assign T_6765 = T_6743[63];
  assign T_6766 = T_6743[65:64];
  assign T_6767 = T_6743[66];
  assign GEN_401 = T_5976 ? T_6717_mie : GEN_372;
  assign GEN_402 = T_5976 ? T_6717_mpie : GEN_373;
  assign T_6796_rocc = T_6822;
  assign T_6796_meip = T_6821;
  assign T_6796_heip = T_6820;
  assign T_6796_seip = T_6819;
  assign T_6796_ueip = T_6818;
  assign T_6796_mtip = T_6817;
  assign T_6796_htip = T_6816;
  assign T_6796_stip = T_6815;
  assign T_6796_utip = T_6814;
  assign T_6796_msip = T_6813;
  assign T_6796_hsip = T_6812;
  assign T_6796_ssip = T_6811;
  assign T_6796_usip = T_6810;
  assign T_6810 = wdata[0];
  assign T_6811 = wdata[1];
  assign T_6812 = wdata[2];
  assign T_6813 = wdata[3];
  assign T_6814 = wdata[4];
  assign T_6815 = wdata[5];
  assign T_6816 = wdata[6];
  assign T_6817 = wdata[7];
  assign T_6818 = wdata[8];
  assign T_6819 = wdata[9];
  assign T_6820 = wdata[10];
  assign T_6821 = wdata[11];
  assign T_6822 = wdata[12];
  assign GEN_11 = {{51'd0}, supported_interrupts};
  assign T_6823 = wdata & GEN_11;
  assign GEN_416 = T_5982 ? T_6823 : reg_mie;
  assign T_6824 = ~ wdata;
  assign T_6826 = T_6824 | 64'h1;
  assign T_6827 = ~ T_6826;
  assign GEN_417 = T_5990 ? T_6827 : {{24'd0}, GEN_347};
  assign GEN_418 = T_5988 ? wdata : reg_mscratch;
  assign T_6828 = wdata[63:2];
  assign GEN_12 = {{2'd0}, T_6828};
  assign T_6829 = GEN_12 << 2;
  assign GEN_419 = T_5978 ? T_6829 : {{32'd0}, reg_mtvec};
  assign T_6831 = wdata & 64'h800000000000001f;
  assign GEN_420 = T_5994 ? T_6831 : GEN_348;
  assign T_6832 = wdata[39:0];
  assign GEN_421 = T_5992 ? T_6832 : GEN_349;
  assign T_6833 = wdata[63:6];
  assign GEN_422 = T_5970 ? wdata : {{57'd0}, T_5579};
  assign GEN_423 = T_5970 ? T_6833 : GEN_39;
  assign GEN_424 = T_5972 ? wdata : {{57'd0}, T_5568};
  assign GEN_425 = T_5972 ? T_6833 : GEN_38;
  assign T_6871_xdebugver = T_6905;
  assign T_6871_ndreset = T_6904;
  assign T_6871_fullreset = T_6903;
  assign T_6871_zero3 = T_6902;
  assign T_6871_ebreakm = T_6901;
  assign T_6871_ebreakh = T_6900;
  assign T_6871_ebreaks = T_6899;
  assign T_6871_ebreaku = T_6822;
  assign T_6871_zero2 = T_6821;
  assign T_6871_stopcycle = T_6820;
  assign T_6871_stoptime = T_6819;
  assign T_6871_cause = T_6894;
  assign T_6871_debugint = T_6815;
  assign T_6871_zero1 = T_6814;
  assign T_6871_halt = T_6813;
  assign T_6871_step = T_6812;
  assign T_6871_prv = T_6889;
  assign T_6889 = wdata[1:0];
  assign T_6894 = wdata[8:6];
  assign T_6899 = wdata[13];
  assign T_6900 = wdata[14];
  assign T_6901 = wdata[15];
  assign T_6902 = wdata[27:16];
  assign T_6903 = wdata[28];
  assign T_6904 = wdata[29];
  assign T_6905 = wdata[31:30];
  assign GEN_443 = T_5998 ? T_6871_halt : reg_dcsr_halt;
  assign GEN_444 = T_5998 ? T_6871_step : reg_dcsr_step;
  assign GEN_445 = T_5998 ? T_6871_ebreakm : reg_dcsr_ebreakm;
  assign GEN_446 = T_6000 ? T_6827 : {{24'd0}, GEN_337};
  assign GEN_447 = T_6002 ? wdata : reg_dscratch;
  assign GEN_17_control_ttype = GEN_42;
  assign GEN_17_control_dmode = GEN_43;
  assign GEN_17_control_maskmax = GEN_44;
  assign GEN_17_control_reserved = GEN_45;
  assign GEN_17_control_action = GEN_46;
  assign GEN_17_control_chain = GEN_47;
  assign GEN_17_control_zero = GEN_48;
  assign GEN_17_control_tmatch = GEN_49;
  assign GEN_17_control_m = GEN_50;
  assign GEN_17_control_h = GEN_51;
  assign GEN_17_control_s = GEN_52;
  assign GEN_17_control_u = GEN_53;
  assign GEN_17_control_x = GEN_54;
  assign GEN_17_control_w = GEN_55;
  assign GEN_17_control_r = GEN_56;
  assign GEN_17_address = GEN_57;
  assign T_6928 = GEN_17_control_dmode == 1'h0;
  assign T_6929 = T_6928 | reg_debug;
  assign T_6962_ttype = T_6992;
  assign T_6962_dmode = T_6991;
  assign T_6962_maskmax = T_6990;
  assign T_6962_reserved = T_6989;
  assign T_6962_action = T_6822;
  assign T_6962_chain = T_6821;
  assign T_6962_zero = T_6986;
  assign T_6962_tmatch = T_6985;
  assign T_6962_m = T_6816;
  assign T_6962_h = T_6815;
  assign T_6962_s = T_6814;
  assign T_6962_u = T_6813;
  assign T_6962_x = T_6812;
  assign T_6962_w = T_6811;
  assign T_6962_r = T_6810;
  assign T_6985 = wdata[8:7];
  assign T_6986 = wdata[10:9];
  assign T_6989 = wdata[52:13];
  assign T_6990 = wdata[58:53];
  assign T_6991 = wdata[59];
  assign T_6992 = wdata[63:60];
  assign T_6993 = T_6962_dmode & reg_debug;
  assign GEN_18 = T_6962_ttype;
  assign GEN_19 = T_6962_dmode;
  assign GEN_467 = 1'h0 == reg_tselect ? GEN_19 : reg_bp_0_control_dmode;
  assign GEN_20 = T_6962_maskmax;
  assign GEN_21 = T_6962_reserved;
  assign GEN_22 = T_6962_action;
  assign GEN_473 = 1'h0 == reg_tselect ? GEN_22 : reg_bp_0_control_action;
  assign GEN_23 = T_6962_chain;
  assign GEN_24 = T_6962_zero;
  assign GEN_25 = T_6962_tmatch;
  assign GEN_479 = 1'h0 == reg_tselect ? GEN_25 : reg_bp_0_control_tmatch;
  assign GEN_26 = T_6962_m;
  assign GEN_27 = T_6962_h;
  assign GEN_28 = T_6962_s;
  assign GEN_29 = T_6962_u;
  assign GEN_30 = T_6962_x;
  assign GEN_489 = 1'h0 == reg_tselect ? GEN_30 : reg_bp_0_control_x;
  assign GEN_31 = T_6962_w;
  assign GEN_491 = 1'h0 == reg_tselect ? GEN_31 : reg_bp_0_control_w;
  assign GEN_32 = T_6962_r;
  assign GEN_493 = 1'h0 == reg_tselect ? GEN_32 : reg_bp_0_control_r;
  assign GEN_33 = T_6993;
  assign GEN_495 = 1'h0 == reg_tselect ? GEN_33 : GEN_467;
  assign T_6994 = T_6993 & T_6962_action;
  assign GEN_34 = T_6994;
  assign GEN_497 = 1'h0 == reg_tselect ? GEN_34 : GEN_473;
  assign GEN_518 = T_5960 ? GEN_495 : reg_bp_0_control_dmode;
  assign GEN_527 = T_5960 ? GEN_497 : reg_bp_0_control_action;
  assign GEN_536 = T_5960 ? GEN_479 : reg_bp_0_control_tmatch;
  assign GEN_551 = T_5960 ? GEN_489 : reg_bp_0_control_x;
  assign GEN_554 = T_5960 ? GEN_491 : reg_bp_0_control_w;
  assign GEN_557 = T_5960 ? GEN_493 : reg_bp_0_control_r;
  assign GEN_35 = wdata[38:0];
  assign GEN_561 = 1'h0 == reg_tselect ? GEN_35 : reg_bp_0_address;
  assign GEN_564 = T_5962 ? GEN_561 : reg_bp_0_address;
  assign GEN_585 = T_6929 ? GEN_518 : reg_bp_0_control_dmode;
  assign GEN_594 = T_6929 ? GEN_527 : reg_bp_0_control_action;
  assign GEN_603 = T_6929 ? GEN_536 : reg_bp_0_control_tmatch;
  assign GEN_618 = T_6929 ? GEN_551 : reg_bp_0_control_x;
  assign GEN_621 = T_6929 ? GEN_554 : reg_bp_0_control_w;
  assign GEN_624 = T_6929 ? GEN_557 : reg_bp_0_control_r;
  assign GEN_629 = T_6929 ? GEN_564 : reg_bp_0_address;
  assign GEN_656 = wen ? GEN_401 : GEN_372;
  assign GEN_657 = wen ? GEN_402 : GEN_373;
  assign GEN_671 = wen ? GEN_416 : reg_mie;
  assign GEN_672 = wen ? GEN_417 : {{24'd0}, GEN_347};
  assign GEN_673 = wen ? GEN_418 : reg_mscratch;
  assign GEN_674 = wen ? GEN_419 : {{32'd0}, reg_mtvec};
  assign GEN_675 = wen ? GEN_420 : GEN_348;
  assign GEN_676 = wen ? GEN_421 : GEN_349;
  assign GEN_677 = wen ? GEN_422 : {{57'd0}, T_5579};
  assign GEN_678 = wen ? GEN_423 : GEN_39;
  assign GEN_679 = wen ? GEN_424 : {{57'd0}, T_5568};
  assign GEN_680 = wen ? GEN_425 : GEN_38;
  assign GEN_698 = wen ? GEN_443 : reg_dcsr_halt;
  assign GEN_699 = wen ? GEN_444 : reg_dcsr_step;
  assign GEN_700 = wen ? GEN_445 : reg_dcsr_ebreakm;
  assign GEN_701 = wen ? GEN_446 : {{24'd0}, GEN_337};
  assign GEN_702 = wen ? GEN_447 : reg_dscratch;
  assign GEN_739 = wen ? GEN_585 : reg_bp_0_control_dmode;
  assign GEN_748 = wen ? GEN_594 : reg_bp_0_control_action;
  assign GEN_757 = wen ? GEN_603 : reg_bp_0_control_tmatch;
  assign GEN_772 = wen ? GEN_618 : reg_bp_0_control_x;
  assign GEN_775 = wen ? GEN_621 : reg_bp_0_control_w;
  assign GEN_778 = wen ? GEN_624 : reg_bp_0_control_r;
  assign GEN_783 = wen ? GEN_629 : reg_bp_0_address;
  assign GEN_785 = reset ? 1'h0 : GEN_748;
  assign GEN_786 = reset ? 1'h0 : GEN_739;
  assign GEN_787 = reset ? 1'h0 : GEN_778;
  assign GEN_788 = reset ? 1'h0 : GEN_775;
  assign GEN_789 = reset ? 1'h0 : GEN_772;
  assign T_7061_control_ttype = T_7096;
  assign T_7061_control_dmode = T_7095;
  assign T_7061_control_maskmax = T_7094;
  assign T_7061_control_reserved = T_7093;
  assign T_7061_control_action = T_7092;
  assign T_7061_control_chain = T_7091;
  assign T_7061_control_zero = T_7090;
  assign T_7061_control_tmatch = T_7089;
  assign T_7061_control_m = T_7088;
  assign T_7061_control_h = T_7087;
  assign T_7061_control_s = T_7086;
  assign T_7061_control_u = T_7085;
  assign T_7061_control_x = T_7084;
  assign T_7061_control_w = T_7083;
  assign T_7061_control_r = T_7082;
  assign T_7061_address = T_7081;
  assign T_7080 = 103'h0;
  assign T_7081 = T_7080[38:0];
  assign T_7082 = T_7080[39];
  assign T_7083 = T_7080[40];
  assign T_7084 = T_7080[41];
  assign T_7085 = T_7080[42];
  assign T_7086 = T_7080[43];
  assign T_7087 = T_7080[44];
  assign T_7088 = T_7080[45];
  assign T_7089 = T_7080[47:46];
  assign T_7090 = T_7080[49:48];
  assign T_7091 = T_7080[50];
  assign T_7092 = T_7080[51];
  assign T_7093 = T_7080[91:52];
  assign T_7094 = T_7080[97:92];
  assign T_7095 = T_7080[98];
  assign T_7096 = T_7080[102:99];
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_13 = GEN_235[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_14 = GEN_236[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_15 = GEN_237[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_16 = GEN_238[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_17 = GEN_239[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_58 = GEN_240[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_59 = GEN_241[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_60 = GEN_242[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_61 = GEN_243[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_62 = GEN_244[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_63 = GEN_245[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_64 = GEN_246[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_65 = GEN_247[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_66 = GEN_248[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_67 = GEN_249[30:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_68 = GEN_250[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_69 = GEN_251[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_70 = GEN_252[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_71 = GEN_253[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_72 = GEN_254[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_73 = GEN_255[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_74 = GEN_256[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_75 = GEN_257[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_76 = GEN_258[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_77 = GEN_259[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_78 = GEN_260[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_79 = GEN_261[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_80 = GEN_262[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_81 = GEN_263[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_82 = GEN_264[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_83 = GEN_265[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_84 = GEN_266[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_85 = GEN_267[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_86 = GEN_268[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_87 = GEN_269[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_88 = GEN_270[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_89 = GEN_271[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_90 = GEN_272[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_91 = GEN_273[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_92 = GEN_274[39:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_93 = GEN_275[5:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_94 = GEN_276[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_95 = GEN_277[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_96 = GEN_278[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_97 = GEN_279[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_98 = GEN_280[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_99 = GEN_281[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_100 = GEN_282[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_101 = GEN_283[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_102 = GEN_284[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_103 = GEN_285[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_104 = GEN_286[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_105 = GEN_287[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_106 = GEN_288[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_107 = GEN_289[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_108 = GEN_290[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_109 = GEN_291[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_110 = GEN_292[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_111 = GEN_293[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_112 = GEN_294[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_113 = GEN_295[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_114 = GEN_296[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_115 = GEN_297[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_116 = GEN_298[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_117 = GEN_299[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_118 = GEN_300[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_119 = GEN_301[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  reg_mstatus_debug = GEN_120[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_121 = {1{$random}};
  reg_mstatus_prv = GEN_121[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_122 = {1{$random}};
  reg_mstatus_sd = GEN_122[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_123 = {1{$random}};
  reg_mstatus_zero3 = GEN_123[30:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_124 = {1{$random}};
  reg_mstatus_sd_rv32 = GEN_124[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_125 = {1{$random}};
  reg_mstatus_zero2 = GEN_125[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_126 = {1{$random}};
  reg_mstatus_vm = GEN_126[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_127 = {1{$random}};
  reg_mstatus_zero1 = GEN_127[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_128 = {1{$random}};
  reg_mstatus_mxr = GEN_128[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_129 = {1{$random}};
  reg_mstatus_pum = GEN_129[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_130 = {1{$random}};
  reg_mstatus_mprv = GEN_130[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_131 = {1{$random}};
  reg_mstatus_xs = GEN_131[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_132 = {1{$random}};
  reg_mstatus_fs = GEN_132[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_133 = {1{$random}};
  reg_mstatus_mpp = GEN_133[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_134 = {1{$random}};
  reg_mstatus_hpp = GEN_134[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_135 = {1{$random}};
  reg_mstatus_spp = GEN_135[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_136 = {1{$random}};
  reg_mstatus_mpie = GEN_136[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_137 = {1{$random}};
  reg_mstatus_hpie = GEN_137[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_138 = {1{$random}};
  reg_mstatus_spie = GEN_138[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_139 = {1{$random}};
  reg_mstatus_upie = GEN_139[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_140 = {1{$random}};
  reg_mstatus_mie = GEN_140[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_141 = {1{$random}};
  reg_mstatus_hie = GEN_141[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_142 = {1{$random}};
  reg_mstatus_sie = GEN_142[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_143 = {1{$random}};
  reg_mstatus_uie = GEN_143[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_144 = {1{$random}};
  reg_dcsr_xdebugver = GEN_144[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_145 = {1{$random}};
  reg_dcsr_ndreset = GEN_145[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_146 = {1{$random}};
  reg_dcsr_fullreset = GEN_146[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_147 = {1{$random}};
  reg_dcsr_zero3 = GEN_147[11:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_148 = {1{$random}};
  reg_dcsr_ebreakm = GEN_148[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_149 = {1{$random}};
  reg_dcsr_ebreakh = GEN_149[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_150 = {1{$random}};
  reg_dcsr_ebreaks = GEN_150[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_151 = {1{$random}};
  reg_dcsr_ebreaku = GEN_151[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_152 = {1{$random}};
  reg_dcsr_zero2 = GEN_152[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_153 = {1{$random}};
  reg_dcsr_stopcycle = GEN_153[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_154 = {1{$random}};
  reg_dcsr_stoptime = GEN_154[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_155 = {1{$random}};
  reg_dcsr_cause = GEN_155[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_156 = {1{$random}};
  reg_dcsr_debugint = GEN_156[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_157 = {1{$random}};
  reg_dcsr_zero1 = GEN_157[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_158 = {1{$random}};
  reg_dcsr_halt = GEN_158[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_159 = {1{$random}};
  reg_dcsr_step = GEN_159[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_160 = {1{$random}};
  reg_dcsr_prv = GEN_160[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_161 = {1{$random}};
  reg_debug = GEN_161[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_162 = {2{$random}};
  reg_dpc = GEN_162[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_163 = {2{$random}};
  reg_dscratch = GEN_163[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_164 = {1{$random}};
  reg_singleStepped = GEN_164[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_165 = {1{$random}};
  reg_tselect = GEN_165[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_166 = {1{$random}};
  reg_bp_0_control_ttype = GEN_166[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_167 = {1{$random}};
  reg_bp_0_control_dmode = GEN_167[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_168 = {1{$random}};
  reg_bp_0_control_maskmax = GEN_168[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_169 = {2{$random}};
  reg_bp_0_control_reserved = GEN_169[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_170 = {1{$random}};
  reg_bp_0_control_action = GEN_170[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_171 = {1{$random}};
  reg_bp_0_control_chain = GEN_171[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_172 = {1{$random}};
  reg_bp_0_control_zero = GEN_172[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_173 = {1{$random}};
  reg_bp_0_control_tmatch = GEN_173[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_174 = {1{$random}};
  reg_bp_0_control_m = GEN_174[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_175 = {1{$random}};
  reg_bp_0_control_h = GEN_175[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_176 = {1{$random}};
  reg_bp_0_control_s = GEN_176[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_177 = {1{$random}};
  reg_bp_0_control_u = GEN_177[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_178 = {1{$random}};
  reg_bp_0_control_x = GEN_178[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_179 = {1{$random}};
  reg_bp_0_control_w = GEN_179[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_180 = {1{$random}};
  reg_bp_0_control_r = GEN_180[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_181 = {2{$random}};
  reg_bp_0_address = GEN_181[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_182 = {1{$random}};
  reg_bp_1_control_ttype = GEN_182[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_183 = {1{$random}};
  reg_bp_1_control_dmode = GEN_183[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_184 = {1{$random}};
  reg_bp_1_control_maskmax = GEN_184[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_185 = {2{$random}};
  reg_bp_1_control_reserved = GEN_185[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_186 = {1{$random}};
  reg_bp_1_control_action = GEN_186[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_187 = {1{$random}};
  reg_bp_1_control_chain = GEN_187[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_188 = {1{$random}};
  reg_bp_1_control_zero = GEN_188[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_189 = {1{$random}};
  reg_bp_1_control_tmatch = GEN_189[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_190 = {1{$random}};
  reg_bp_1_control_m = GEN_190[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_191 = {1{$random}};
  reg_bp_1_control_h = GEN_191[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_192 = {1{$random}};
  reg_bp_1_control_s = GEN_192[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_193 = {1{$random}};
  reg_bp_1_control_u = GEN_193[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_194 = {1{$random}};
  reg_bp_1_control_x = GEN_194[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_195 = {1{$random}};
  reg_bp_1_control_w = GEN_195[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_196 = {1{$random}};
  reg_bp_1_control_r = GEN_196[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_197 = {2{$random}};
  reg_bp_1_address = GEN_197[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_198 = {2{$random}};
  reg_mie = GEN_198[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_199 = {2{$random}};
  reg_mideleg = GEN_199[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_200 = {2{$random}};
  reg_medeleg = GEN_200[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_201 = {1{$random}};
  reg_mip_rocc = GEN_201[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_202 = {1{$random}};
  reg_mip_meip = GEN_202[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_203 = {1{$random}};
  reg_mip_heip = GEN_203[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_204 = {1{$random}};
  reg_mip_seip = GEN_204[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_205 = {1{$random}};
  reg_mip_ueip = GEN_205[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_206 = {1{$random}};
  reg_mip_mtip = GEN_206[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_207 = {1{$random}};
  reg_mip_htip = GEN_207[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_208 = {1{$random}};
  reg_mip_stip = GEN_208[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_209 = {1{$random}};
  reg_mip_utip = GEN_209[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_210 = {1{$random}};
  reg_mip_msip = GEN_210[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_211 = {1{$random}};
  reg_mip_hsip = GEN_211[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_212 = {1{$random}};
  reg_mip_ssip = GEN_212[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_213 = {1{$random}};
  reg_mip_usip = GEN_213[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_214 = {2{$random}};
  reg_mepc = GEN_214[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_215 = {2{$random}};
  reg_mcause = GEN_215[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_216 = {2{$random}};
  reg_mbadaddr = GEN_216[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_217 = {2{$random}};
  reg_mscratch = GEN_217[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_218 = {1{$random}};
  reg_mtvec = GEN_218[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_219 = {1{$random}};
  reg_mucounteren = GEN_219[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_220 = {1{$random}};
  reg_mscounteren = GEN_220[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_221 = {2{$random}};
  reg_sepc = GEN_221[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_222 = {2{$random}};
  reg_scause = GEN_222[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_223 = {2{$random}};
  reg_sbadaddr = GEN_223[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_224 = {2{$random}};
  reg_sscratch = GEN_224[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_225 = {2{$random}};
  reg_stvec = GEN_225[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_226 = {1{$random}};
  reg_sptbr_asid = GEN_226[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_227 = {2{$random}};
  reg_sptbr_ppn = GEN_227[37:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_228 = {1{$random}};
  reg_wfi = GEN_228[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_229 = {1{$random}};
  reg_fflags = GEN_229[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_230 = {1{$random}};
  reg_frm = GEN_230[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_231 = {1{$random}};
  T_5567 = GEN_231[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_232 = {2{$random}};
  T_5570 = GEN_232[57:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_233 = {1{$random}};
  T_5578 = GEN_233[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_234 = {2{$random}};
  T_5581 = GEN_234[57:0];
  `endif
  GEN_235 = {1{$random}};
  GEN_236 = {1{$random}};
  GEN_237 = {1{$random}};
  GEN_238 = {1{$random}};
  GEN_239 = {1{$random}};
  GEN_240 = {1{$random}};
  GEN_241 = {1{$random}};
  GEN_242 = {1{$random}};
  GEN_243 = {1{$random}};
  GEN_244 = {2{$random}};
  GEN_245 = {2{$random}};
  GEN_246 = {1{$random}};
  GEN_247 = {1{$random}};
  GEN_248 = {1{$random}};
  GEN_249 = {1{$random}};
  GEN_250 = {1{$random}};
  GEN_251 = {1{$random}};
  GEN_252 = {1{$random}};
  GEN_253 = {1{$random}};
  GEN_254 = {1{$random}};
  GEN_255 = {1{$random}};
  GEN_256 = {1{$random}};
  GEN_257 = {1{$random}};
  GEN_258 = {1{$random}};
  GEN_259 = {1{$random}};
  GEN_260 = {1{$random}};
  GEN_261 = {1{$random}};
  GEN_262 = {1{$random}};
  GEN_263 = {1{$random}};
  GEN_264 = {1{$random}};
  GEN_265 = {1{$random}};
  GEN_266 = {1{$random}};
  GEN_267 = {1{$random}};
  GEN_268 = {1{$random}};
  GEN_269 = {1{$random}};
  GEN_270 = {1{$random}};
  GEN_271 = {1{$random}};
  GEN_272 = {1{$random}};
  GEN_273 = {1{$random}};
  GEN_274 = {2{$random}};
  GEN_275 = {1{$random}};
  GEN_276 = {1{$random}};
  GEN_277 = {1{$random}};
  GEN_278 = {2{$random}};
  GEN_279 = {1{$random}};
  GEN_280 = {1{$random}};
  GEN_281 = {2{$random}};
  GEN_282 = {2{$random}};
  GEN_283 = {1{$random}};
  GEN_284 = {1{$random}};
  GEN_285 = {1{$random}};
  GEN_286 = {1{$random}};
  GEN_287 = {1{$random}};
  GEN_288 = {1{$random}};
  GEN_289 = {1{$random}};
  GEN_290 = {1{$random}};
  GEN_291 = {1{$random}};
  GEN_292 = {1{$random}};
  GEN_293 = {1{$random}};
  GEN_294 = {1{$random}};
  GEN_295 = {1{$random}};
  GEN_296 = {2{$random}};
  GEN_297 = {1{$random}};
  GEN_298 = {1{$random}};
  GEN_299 = {3{$random}};
  GEN_300 = {1{$random}};
  GEN_301 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      reg_mstatus_debug <= reset_mstatus_debug;
    end
    if(reset) begin
      reg_mstatus_prv <= reset_mstatus_prv;
    end else begin
      reg_mstatus_prv <= 2'h3;
    end
    if(reset) begin
      reg_mstatus_sd <= reset_mstatus_sd;
    end
    if(reset) begin
      reg_mstatus_zero3 <= reset_mstatus_zero3;
    end
    if(reset) begin
      reg_mstatus_sd_rv32 <= reset_mstatus_sd_rv32;
    end
    if(reset) begin
      reg_mstatus_zero2 <= reset_mstatus_zero2;
    end
    if(reset) begin
      reg_mstatus_vm <= reset_mstatus_vm;
    end
    if(reset) begin
      reg_mstatus_zero1 <= reset_mstatus_zero1;
    end
    if(reset) begin
      reg_mstatus_mxr <= reset_mstatus_mxr;
    end
    if(reset) begin
      reg_mstatus_pum <= reset_mstatus_pum;
    end
    if(reset) begin
      reg_mstatus_mprv <= reset_mstatus_mprv;
    end
    if(reset) begin
      reg_mstatus_xs <= reset_mstatus_xs;
    end
    if(reset) begin
      reg_mstatus_fs <= reset_mstatus_fs;
    end
    if(reset) begin
      reg_mstatus_mpp <= reset_mstatus_mpp;
    end else begin
      if(insn_ret) begin
        if(T_6220) begin
          reg_mstatus_mpp <= 2'h3;
        end else begin
          if(exception) begin
            if(T_6376) begin
              reg_mstatus_mpp <= 2'h3;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6376) begin
            reg_mstatus_mpp <= 2'h3;
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_hpp <= reset_mstatus_hpp;
    end
    if(reset) begin
      reg_mstatus_spp <= reset_mstatus_spp;
    end else begin
      reg_mstatus_spp <= GEN_344[0];
    end
    if(reset) begin
      reg_mstatus_mpie <= reset_mstatus_mpie;
    end else begin
      if(wen) begin
        if(T_5976) begin
          reg_mstatus_mpie <= T_6717_mpie;
        end else begin
          if(insn_ret) begin
            if(T_6220) begin
              reg_mstatus_mpie <= 1'h0;
            end else begin
              if(exception) begin
                if(T_6376) begin
                  reg_mstatus_mpie <= T_6345;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6376) begin
                reg_mstatus_mpie <= T_6345;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6220) begin
            reg_mstatus_mpie <= 1'h0;
          end else begin
            if(exception) begin
              if(T_6376) begin
                reg_mstatus_mpie <= T_6345;
              end
            end
          end
        end else begin
          if(exception) begin
            if(T_6376) begin
              reg_mstatus_mpie <= T_6345;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_hpie <= reset_mstatus_hpie;
    end
    if(reset) begin
      reg_mstatus_spie <= reset_mstatus_spie;
    end
    if(reset) begin
      reg_mstatus_upie <= reset_mstatus_upie;
    end
    if(reset) begin
      reg_mstatus_mie <= reset_mstatus_mie;
    end else begin
      if(wen) begin
        if(T_5976) begin
          reg_mstatus_mie <= T_6717_mie;
        end else begin
          if(insn_ret) begin
            if(T_6220) begin
              if(T_6405) begin
                reg_mstatus_mie <= reg_mstatus_mpie;
              end else begin
                if(exception) begin
                  if(T_6376) begin
                    reg_mstatus_mie <= 1'h0;
                  end
                end
              end
            end else begin
              if(exception) begin
                if(T_6376) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6376) begin
                reg_mstatus_mie <= 1'h0;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6220) begin
            if(T_6405) begin
              reg_mstatus_mie <= reg_mstatus_mpie;
            end else begin
              if(exception) begin
                if(T_6376) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            reg_mstatus_mie <= GEN_352;
          end
        end else begin
          reg_mstatus_mie <= GEN_352;
        end
      end
    end
    if(reset) begin
      reg_mstatus_hie <= reset_mstatus_hie;
    end
    if(reset) begin
      reg_mstatus_sie <= reset_mstatus_sie;
    end
    if(reset) begin
      reg_mstatus_uie <= reset_mstatus_uie;
    end
    if(reset) begin
      reg_dcsr_xdebugver <= reset_dcsr_xdebugver;
    end
    if(reset) begin
      reg_dcsr_ndreset <= reset_dcsr_ndreset;
    end
    if(reset) begin
      reg_dcsr_fullreset <= reset_dcsr_fullreset;
    end
    if(reset) begin
      reg_dcsr_zero3 <= reset_dcsr_zero3;
    end
    if(reset) begin
      reg_dcsr_ebreakm <= reset_dcsr_ebreakm;
    end else begin
      if(wen) begin
        if(T_5998) begin
          reg_dcsr_ebreakm <= T_6871_ebreakm;
        end
      end
    end
    if(reset) begin
      reg_dcsr_ebreakh <= reset_dcsr_ebreakh;
    end
    if(reset) begin
      reg_dcsr_ebreaks <= reset_dcsr_ebreaks;
    end
    if(reset) begin
      reg_dcsr_ebreaku <= reset_dcsr_ebreaku;
    end
    if(reset) begin
      reg_dcsr_zero2 <= reset_dcsr_zero2;
    end
    if(reset) begin
      reg_dcsr_stopcycle <= reset_dcsr_stopcycle;
    end
    if(reset) begin
      reg_dcsr_stoptime <= reset_dcsr_stoptime;
    end
    if(reset) begin
      reg_dcsr_cause <= reset_dcsr_cause;
    end else begin
      if(exception) begin
        if(T_6307) begin
          if(reg_singleStepped) begin
            reg_dcsr_cause <= 3'h4;
          end else begin
            reg_dcsr_cause <= {{1'd0}, T_6372};
          end
        end
      end
    end
    if(reset) begin
      reg_dcsr_debugint <= reset_dcsr_debugint;
    end else begin
      reg_dcsr_debugint <= io_prci_interrupts_debug;
    end
    if(reset) begin
      reg_dcsr_zero1 <= reset_dcsr_zero1;
    end
    if(reset) begin
      reg_dcsr_halt <= reset_dcsr_halt;
    end else begin
      if(wen) begin
        if(T_5998) begin
          reg_dcsr_halt <= T_6871_halt;
        end
      end
    end
    if(reset) begin
      reg_dcsr_step <= reset_dcsr_step;
    end else begin
      if(wen) begin
        if(T_5998) begin
          reg_dcsr_step <= T_6871_step;
        end
      end
    end
    if(reset) begin
      reg_dcsr_prv <= reset_dcsr_prv;
    end else begin
      if(exception) begin
        if(T_6307) begin
          reg_dcsr_prv <= 2'h3;
        end
      end
    end
    if(reset) begin
      reg_debug <= 1'h0;
    end else begin
      if(insn_ret) begin
        if(T_6218) begin
          reg_debug <= 1'h0;
        end else begin
          if(exception) begin
            if(T_6307) begin
              reg_debug <= 1'h1;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6307) begin
            reg_debug <= 1'h1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_dpc <= GEN_701[39:0];
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6002) begin
          reg_dscratch <= wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5320) begin
        reg_singleStepped <= 1'h0;
      end else begin
        if(T_5317) begin
          reg_singleStepped <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_tselect <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_ttype <= 4'h2;
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_dmode <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6929) begin
            if(T_5960) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_dmode <= GEN_33;
              end else begin
                if(1'h0 == reg_tselect) begin
                  reg_bp_0_control_dmode <= GEN_19;
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_maskmax <= 6'h4;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_reserved <= 40'h0;
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_action <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6929) begin
            if(T_5960) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_action <= GEN_34;
              end else begin
                if(1'h0 == reg_tselect) begin
                  reg_bp_0_control_action <= GEN_22;
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_chain <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_zero <= 2'h0;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6929) begin
          if(T_5960) begin
            if(1'h0 == reg_tselect) begin
              reg_bp_0_control_tmatch <= GEN_25;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_m <= 1'h1;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_h <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_s <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_u <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_x <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6929) begin
            if(T_5960) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_x <= GEN_30;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_w <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6929) begin
            if(T_5960) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_w <= GEN_31;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_r <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6929) begin
            if(T_5960) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_r <= GEN_32;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6929) begin
          if(T_5962) begin
            if(1'h0 == reg_tselect) begin
              reg_bp_0_address <= GEN_35;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_ttype <= T_7061_control_ttype;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_dmode <= T_7061_control_dmode;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_maskmax <= T_7061_control_maskmax;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_reserved <= T_7061_control_reserved;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_action <= T_7061_control_action;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_chain <= T_7061_control_chain;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_zero <= T_7061_control_zero;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_tmatch <= T_7061_control_tmatch;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_m <= T_7061_control_m;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_h <= T_7061_control_h;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_s <= T_7061_control_s;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_u <= T_7061_control_u;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_x <= T_7061_control_x;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_w <= T_7061_control_w;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_r <= T_7061_control_r;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_address <= T_7061_address;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5982) begin
          reg_mie <= T_6823;
        end
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_meip <= io_prci_interrupts_meip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_seip <= io_prci_interrupts_seip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_mtip <= io_prci_interrupts_mtip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_msip <= io_prci_interrupts_msip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mepc <= GEN_672[39:0];
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5994) begin
          reg_mcause <= T_6831;
        end else begin
          if(exception) begin
            if(T_6376) begin
              if(T_6278) begin
                reg_mcause <= io_cause;
              end else begin
                reg_mcause <= {{60'd0}, T_6285};
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6376) begin
            if(T_6278) begin
              reg_mcause <= io_cause;
            end else begin
              reg_mcause <= {{60'd0}, T_6285};
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5992) begin
          reg_mbadaddr <= T_6832;
        end else begin
          if(exception) begin
            if(T_6376) begin
              if(T_6365) begin
                reg_mbadaddr <= io_badaddr;
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6376) begin
            if(T_6365) begin
              reg_mbadaddr <= io_badaddr;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5988) begin
          reg_mscratch <= wdata;
        end
      end
    end
    if(reset) begin
      reg_mtvec <= 32'h1010;
    end else begin
      reg_mtvec <= GEN_674[31:0];
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_sptbr_asid <= 7'h0;
    end
    if(1'h0) begin
    end
    if(reset) begin
      reg_wfi <= 1'h0;
    end else begin
      if(T_6275) begin
        reg_wfi <= 1'h0;
      end else begin
        if(insn_wfi) begin
          reg_wfi <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_fcsr_flags_valid) begin
        reg_fflags <= T_6666;
      end
    end
    if(1'h0) begin
    end
    if(reset) begin
      T_5567 <= 6'h0;
    end else begin
      T_5567 <= GEN_679[5:0];
    end
    if(reset) begin
      T_5570 <= 58'h0;
    end else begin
      if(wen) begin
        if(T_5972) begin
          T_5570 <= T_6833;
        end else begin
          if(T_5571) begin
            T_5570 <= T_5574;
          end
        end
      end else begin
        if(T_5571) begin
          T_5570 <= T_5574;
        end
      end
    end
    if(reset) begin
      T_5578 <= 6'h0;
    end else begin
      T_5578 <= GEN_677[5:0];
    end
    if(reset) begin
      T_5581 <= 58'h0;
    end else begin
      if(wen) begin
        if(T_5970) begin
          T_5581 <= T_6833;
        end else begin
          if(T_5582) begin
            T_5581 <= T_5585;
          end
        end
      end else begin
        if(T_5582) begin
          T_5581 <= T_5585;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at csr.scala:204 assert(!io.singleStep || io.retire <= UInt(1))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_5337) begin
          $fwrite(32'h80000002,"Assertion failed\n    at csr.scala:205 assert(!reg_singleStepped || io.retire === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_5337) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_6421) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at csr.scala:478 assert(PopCount(insn_ret :: io.exception :: io.csr_xcpt :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_6421) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BreakpointUnit(
  input   clk,
  input   reset,
  input   io_status_debug,
  input  [1:0] io_status_prv,
  input   io_status_sd,
  input  [30:0] io_status_zero3,
  input   io_status_sd_rv32,
  input  [1:0] io_status_zero2,
  input  [4:0] io_status_vm,
  input  [3:0] io_status_zero1,
  input   io_status_mxr,
  input   io_status_pum,
  input   io_status_mprv,
  input  [1:0] io_status_xs,
  input  [1:0] io_status_fs,
  input  [1:0] io_status_mpp,
  input  [1:0] io_status_hpp,
  input   io_status_spp,
  input   io_status_mpie,
  input   io_status_hpie,
  input   io_status_spie,
  input   io_status_upie,
  input   io_status_mie,
  input   io_status_hie,
  input   io_status_sie,
  input   io_status_uie,
  input  [3:0] io_bp_0_control_ttype,
  input   io_bp_0_control_dmode,
  input  [5:0] io_bp_0_control_maskmax,
  input  [39:0] io_bp_0_control_reserved,
  input   io_bp_0_control_action,
  input   io_bp_0_control_chain,
  input  [1:0] io_bp_0_control_zero,
  input  [1:0] io_bp_0_control_tmatch,
  input   io_bp_0_control_m,
  input   io_bp_0_control_h,
  input   io_bp_0_control_s,
  input   io_bp_0_control_u,
  input   io_bp_0_control_x,
  input   io_bp_0_control_w,
  input   io_bp_0_control_r,
  input  [38:0] io_bp_0_address,
  input  [38:0] io_pc,
  input  [38:0] io_ea,
  output  io_xcpt_if,
  output  io_xcpt_ld,
  output  io_xcpt_st,
  output  io_debug_if,
  output  io_debug_ld,
  output  io_debug_st
);
  wire  T_212;
  wire [1:0] T_213;
  wire [1:0] T_214;
  wire [3:0] T_215;
  wire [3:0] T_216;
  wire  T_217;
  wire  T_218;
  wire  T_220;
  wire  T_221;
  wire  T_222;
  wire  T_223;
  wire  T_224;
  wire [38:0] T_225;
  wire  T_227;
  wire  T_228;
  wire  T_229;
  wire  T_230;
  wire  T_231;
  wire  T_232;
  wire [1:0] T_233;
  wire [1:0] T_234;
  wire [3:0] T_235;
  wire [38:0] GEN_6;
  wire [38:0] T_236;
  wire [38:0] T_237;
  wire [38:0] T_248;
  wire  T_249;
  wire  T_250;
  wire  T_251;
  wire  T_253;
  wire  T_284;
  wire  T_286;
  wire  T_288;
  wire  T_290;
  wire [38:0] T_291;
  wire [38:0] T_302;
  wire  T_315;
  wire  T_316;
  wire  T_317;
  wire  T_319;
  wire  T_320;
  wire  T_322;
  wire  GEN_0;
  wire  GEN_1;
  wire  T_323;
  wire  GEN_2;
  wire  GEN_3;
  wire  T_326;
  wire  GEN_4;
  wire  GEN_5;
  assign io_xcpt_if = GEN_4;
  assign io_xcpt_ld = GEN_0;
  assign io_xcpt_st = GEN_2;
  assign io_debug_if = GEN_5;
  assign io_debug_ld = GEN_1;
  assign io_debug_st = GEN_3;
  assign T_212 = io_status_debug == 1'h0;
  assign T_213 = {io_bp_0_control_s,io_bp_0_control_u};
  assign T_214 = {io_bp_0_control_m,io_bp_0_control_h};
  assign T_215 = {T_214,T_213};
  assign T_216 = T_215 >> io_status_prv;
  assign T_217 = T_216[0];
  assign T_218 = T_212 & T_217;
  assign T_220 = T_218 & io_bp_0_control_r;
  assign T_221 = io_bp_0_control_tmatch[1];
  assign T_222 = io_ea >= io_bp_0_address;
  assign T_223 = io_bp_0_control_tmatch[0];
  assign T_224 = T_222 ^ T_223;
  assign T_225 = ~ io_ea;
  assign T_227 = io_bp_0_address[0];
  assign T_228 = T_223 & T_227;
  assign T_229 = io_bp_0_address[1];
  assign T_230 = T_228 & T_229;
  assign T_231 = io_bp_0_address[2];
  assign T_232 = T_230 & T_231;
  assign T_233 = {T_228,T_223};
  assign T_234 = {T_232,T_230};
  assign T_235 = {T_234,T_233};
  assign GEN_6 = {{35'd0}, T_235};
  assign T_236 = T_225 | GEN_6;
  assign T_237 = ~ io_bp_0_address;
  assign T_248 = T_237 | GEN_6;
  assign T_249 = T_236 == T_248;
  assign T_250 = T_221 ? T_224 : T_249;
  assign T_251 = T_220 & T_250;
  assign T_253 = T_218 & io_bp_0_control_w;
  assign T_284 = T_253 & T_250;
  assign T_286 = T_218 & io_bp_0_control_x;
  assign T_288 = io_pc >= io_bp_0_address;
  assign T_290 = T_288 ^ T_223;
  assign T_291 = ~ io_pc;
  assign T_302 = T_291 | GEN_6;
  assign T_315 = T_302 == T_248;
  assign T_316 = T_221 ? T_290 : T_315;
  assign T_317 = T_286 & T_316;
  assign T_319 = io_bp_0_control_chain == 1'h0;
  assign T_320 = T_319 & T_251;
  assign T_322 = io_bp_0_control_action == 1'h0;
  assign GEN_0 = T_320 ? T_322 : 1'h0;
  assign GEN_1 = T_320 ? io_bp_0_control_action : 1'h0;
  assign T_323 = T_319 & T_284;
  assign GEN_2 = T_323 ? T_322 : 1'h0;
  assign GEN_3 = T_323 ? io_bp_0_control_action : 1'h0;
  assign T_326 = T_319 & T_317;
  assign GEN_4 = T_326 ? T_322 : 1'h0;
  assign GEN_5 = T_326 ? io_bp_0_control_action : 1'h0;
endmodule
module ALU(
  input   clk,
  input   reset,
  input   io_dw,
  input  [3:0] io_fn,
  input  [63:0] io_in2,
  input  [63:0] io_in1,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output  io_cmp_out
);
  wire  T_7;
  wire [63:0] T_8;
  wire [63:0] in2_inv;
  wire [63:0] in1_xor_in2;
  wire [64:0] T_9;
  wire [63:0] T_10;
  wire [63:0] GEN_1;
  wire [64:0] T_12;
  wire [63:0] T_13;
  wire  T_14;
  wire  T_17;
  wire  T_19;
  wire  T_20;
  wire  T_21;
  wire  T_22;
  wire  T_23;
  wire  T_24;
  wire  T_27;
  wire  T_28;
  wire  T_29;
  wire  T_30;
  wire  T_32;
  wire  T_33;
  wire [31:0] T_37;
  wire [31:0] T_39;
  wire [31:0] T_40;
  wire  T_41;
  wire  T_43;
  wire [4:0] T_44;
  wire [5:0] shamt;
  wire [31:0] T_45;
  wire [63:0] shin_r;
  wire  T_46;
  wire  T_47;
  wire  T_48;
  wire [31:0] T_53;
  wire [63:0] T_54;
  wire [31:0] T_55;
  wire [63:0] GEN_2;
  wire [63:0] T_56;
  wire [63:0] T_58;
  wire [63:0] T_59;
  wire [47:0] T_63;
  wire [63:0] GEN_3;
  wire [63:0] T_64;
  wire [47:0] T_65;
  wire [63:0] GEN_4;
  wire [63:0] T_66;
  wire [63:0] T_68;
  wire [63:0] T_69;
  wire [55:0] T_73;
  wire [63:0] GEN_5;
  wire [63:0] T_74;
  wire [55:0] T_75;
  wire [63:0] GEN_6;
  wire [63:0] T_76;
  wire [63:0] T_78;
  wire [63:0] T_79;
  wire [59:0] T_83;
  wire [63:0] GEN_7;
  wire [63:0] T_84;
  wire [59:0] T_85;
  wire [63:0] GEN_8;
  wire [63:0] T_86;
  wire [63:0] T_88;
  wire [63:0] T_89;
  wire [61:0] T_93;
  wire [63:0] GEN_9;
  wire [63:0] T_94;
  wire [61:0] T_95;
  wire [63:0] GEN_10;
  wire [63:0] T_96;
  wire [63:0] T_98;
  wire [63:0] T_99;
  wire [62:0] T_103;
  wire [63:0] GEN_11;
  wire [63:0] T_104;
  wire [62:0] T_105;
  wire [63:0] GEN_12;
  wire [63:0] T_106;
  wire [63:0] T_108;
  wire [63:0] T_109;
  wire [63:0] shin;
  wire  T_111;
  wire  T_112;
  wire [64:0] T_113;
  wire [64:0] T_114;
  wire [64:0] T_115;
  wire [63:0] shout_r;
  wire [31:0] T_120;
  wire [63:0] T_121;
  wire [31:0] T_122;
  wire [63:0] GEN_13;
  wire [63:0] T_123;
  wire [63:0] T_125;
  wire [63:0] T_126;
  wire [47:0] T_130;
  wire [63:0] GEN_14;
  wire [63:0] T_131;
  wire [47:0] T_132;
  wire [63:0] GEN_15;
  wire [63:0] T_133;
  wire [63:0] T_135;
  wire [63:0] T_136;
  wire [55:0] T_140;
  wire [63:0] GEN_16;
  wire [63:0] T_141;
  wire [55:0] T_142;
  wire [63:0] GEN_17;
  wire [63:0] T_143;
  wire [63:0] T_145;
  wire [63:0] T_146;
  wire [59:0] T_150;
  wire [63:0] GEN_18;
  wire [63:0] T_151;
  wire [59:0] T_152;
  wire [63:0] GEN_19;
  wire [63:0] T_153;
  wire [63:0] T_155;
  wire [63:0] T_156;
  wire [61:0] T_160;
  wire [63:0] GEN_20;
  wire [63:0] T_161;
  wire [61:0] T_162;
  wire [63:0] GEN_21;
  wire [63:0] T_163;
  wire [63:0] T_165;
  wire [63:0] T_166;
  wire [62:0] T_170;
  wire [63:0] GEN_22;
  wire [63:0] T_171;
  wire [62:0] T_172;
  wire [63:0] GEN_23;
  wire [63:0] T_173;
  wire [63:0] T_175;
  wire [63:0] shout_l;
  wire [63:0] T_180;
  wire  T_181;
  wire [63:0] T_183;
  wire [63:0] shout;
  wire  T_184;
  wire  T_185;
  wire  T_186;
  wire [63:0] T_188;
  wire  T_190;
  wire  T_191;
  wire [63:0] T_192;
  wire [63:0] T_194;
  wire [63:0] logic$;
  wire  T_195;
  wire  T_196;
  wire  T_197;
  wire  T_198;
  wire  T_199;
  wire  T_200;
  wire [63:0] GEN_24;
  wire [63:0] T_201;
  wire [63:0] shift_logic;
  wire  T_202;
  wire  T_203;
  wire  T_204;
  wire [63:0] out;
  wire  T_205;
  wire  T_206;
  wire [31:0] T_210;
  wire [31:0] T_211;
  wire [63:0] T_212;
  wire [63:0] GEN_0;
  assign io_out = GEN_0;
  assign io_adder_out = T_13;
  assign io_cmp_out = T_30;
  assign T_7 = io_fn[3];
  assign T_8 = ~ io_in2;
  assign in2_inv = T_7 ? T_8 : io_in2;
  assign in1_xor_in2 = io_in1 ^ in2_inv;
  assign T_9 = io_in1 + in2_inv;
  assign T_10 = T_9[63:0];
  assign GEN_1 = {{63'd0}, T_7};
  assign T_12 = T_10 + GEN_1;
  assign T_13 = T_12[63:0];
  assign T_14 = io_fn[0];
  assign T_17 = T_7 == 1'h0;
  assign T_19 = in1_xor_in2 == 64'h0;
  assign T_20 = io_in1[63];
  assign T_21 = io_in2[63];
  assign T_22 = T_20 == T_21;
  assign T_23 = io_adder_out[63];
  assign T_24 = io_fn[1];
  assign T_27 = T_24 ? T_21 : T_20;
  assign T_28 = T_22 ? T_23 : T_27;
  assign T_29 = T_17 ? T_19 : T_28;
  assign T_30 = T_14 ^ T_29;
  assign T_32 = io_in1[31];
  assign T_33 = T_7 & T_32;
  assign T_37 = T_33 ? 32'hffffffff : 32'h0;
  assign T_39 = io_in1[63:32];
  assign T_40 = io_dw ? T_39 : T_37;
  assign T_41 = io_in2[5];
  assign T_43 = T_41 & io_dw;
  assign T_44 = io_in2[4:0];
  assign shamt = {T_43,T_44};
  assign T_45 = io_in1[31:0];
  assign shin_r = {T_40,T_45};
  assign T_46 = io_fn == 4'h5;
  assign T_47 = io_fn == 4'hb;
  assign T_48 = T_46 | T_47;
  assign T_53 = shin_r[63:32];
  assign T_54 = {{32'd0}, T_53};
  assign T_55 = shin_r[31:0];
  assign GEN_2 = {{32'd0}, T_55};
  assign T_56 = GEN_2 << 32;
  assign T_58 = T_56 & 64'hffffffff00000000;
  assign T_59 = T_54 | T_58;
  assign T_63 = T_59[63:16];
  assign GEN_3 = {{16'd0}, T_63};
  assign T_64 = GEN_3 & 64'hffff0000ffff;
  assign T_65 = T_59[47:0];
  assign GEN_4 = {{16'd0}, T_65};
  assign T_66 = GEN_4 << 16;
  assign T_68 = T_66 & 64'hffff0000ffff0000;
  assign T_69 = T_64 | T_68;
  assign T_73 = T_69[63:8];
  assign GEN_5 = {{8'd0}, T_73};
  assign T_74 = GEN_5 & 64'hff00ff00ff00ff;
  assign T_75 = T_69[55:0];
  assign GEN_6 = {{8'd0}, T_75};
  assign T_76 = GEN_6 << 8;
  assign T_78 = T_76 & 64'hff00ff00ff00ff00;
  assign T_79 = T_74 | T_78;
  assign T_83 = T_79[63:4];
  assign GEN_7 = {{4'd0}, T_83};
  assign T_84 = GEN_7 & 64'hf0f0f0f0f0f0f0f;
  assign T_85 = T_79[59:0];
  assign GEN_8 = {{4'd0}, T_85};
  assign T_86 = GEN_8 << 4;
  assign T_88 = T_86 & 64'hf0f0f0f0f0f0f0f0;
  assign T_89 = T_84 | T_88;
  assign T_93 = T_89[63:2];
  assign GEN_9 = {{2'd0}, T_93};
  assign T_94 = GEN_9 & 64'h3333333333333333;
  assign T_95 = T_89[61:0];
  assign GEN_10 = {{2'd0}, T_95};
  assign T_96 = GEN_10 << 2;
  assign T_98 = T_96 & 64'hcccccccccccccccc;
  assign T_99 = T_94 | T_98;
  assign T_103 = T_99[63:1];
  assign GEN_11 = {{1'd0}, T_103};
  assign T_104 = GEN_11 & 64'h5555555555555555;
  assign T_105 = T_99[62:0];
  assign GEN_12 = {{1'd0}, T_105};
  assign T_106 = GEN_12 << 1;
  assign T_108 = T_106 & 64'haaaaaaaaaaaaaaaa;
  assign T_109 = T_104 | T_108;
  assign shin = T_48 ? shin_r : T_109;
  assign T_111 = shin[63];
  assign T_112 = T_7 & T_111;
  assign T_113 = {T_112,shin};
  assign T_114 = $signed(T_113);
  assign T_115 = $signed(T_114) >>> shamt;
  assign shout_r = T_115[63:0];
  assign T_120 = shout_r[63:32];
  assign T_121 = {{32'd0}, T_120};
  assign T_122 = shout_r[31:0];
  assign GEN_13 = {{32'd0}, T_122};
  assign T_123 = GEN_13 << 32;
  assign T_125 = T_123 & 64'hffffffff00000000;
  assign T_126 = T_121 | T_125;
  assign T_130 = T_126[63:16];
  assign GEN_14 = {{16'd0}, T_130};
  assign T_131 = GEN_14 & 64'hffff0000ffff;
  assign T_132 = T_126[47:0];
  assign GEN_15 = {{16'd0}, T_132};
  assign T_133 = GEN_15 << 16;
  assign T_135 = T_133 & 64'hffff0000ffff0000;
  assign T_136 = T_131 | T_135;
  assign T_140 = T_136[63:8];
  assign GEN_16 = {{8'd0}, T_140};
  assign T_141 = GEN_16 & 64'hff00ff00ff00ff;
  assign T_142 = T_136[55:0];
  assign GEN_17 = {{8'd0}, T_142};
  assign T_143 = GEN_17 << 8;
  assign T_145 = T_143 & 64'hff00ff00ff00ff00;
  assign T_146 = T_141 | T_145;
  assign T_150 = T_146[63:4];
  assign GEN_18 = {{4'd0}, T_150};
  assign T_151 = GEN_18 & 64'hf0f0f0f0f0f0f0f;
  assign T_152 = T_146[59:0];
  assign GEN_19 = {{4'd0}, T_152};
  assign T_153 = GEN_19 << 4;
  assign T_155 = T_153 & 64'hf0f0f0f0f0f0f0f0;
  assign T_156 = T_151 | T_155;
  assign T_160 = T_156[63:2];
  assign GEN_20 = {{2'd0}, T_160};
  assign T_161 = GEN_20 & 64'h3333333333333333;
  assign T_162 = T_156[61:0];
  assign GEN_21 = {{2'd0}, T_162};
  assign T_163 = GEN_21 << 2;
  assign T_165 = T_163 & 64'hcccccccccccccccc;
  assign T_166 = T_161 | T_165;
  assign T_170 = T_166[63:1];
  assign GEN_22 = {{1'd0}, T_170};
  assign T_171 = GEN_22 & 64'h5555555555555555;
  assign T_172 = T_166[62:0];
  assign GEN_23 = {{1'd0}, T_172};
  assign T_173 = GEN_23 << 1;
  assign T_175 = T_173 & 64'haaaaaaaaaaaaaaaa;
  assign shout_l = T_171 | T_175;
  assign T_180 = T_48 ? shout_r : 64'h0;
  assign T_181 = io_fn == 4'h1;
  assign T_183 = T_181 ? shout_l : 64'h0;
  assign shout = T_180 | T_183;
  assign T_184 = io_fn == 4'h4;
  assign T_185 = io_fn == 4'h6;
  assign T_186 = T_184 | T_185;
  assign T_188 = T_186 ? in1_xor_in2 : 64'h0;
  assign T_190 = io_fn == 4'h7;
  assign T_191 = T_185 | T_190;
  assign T_192 = io_in1 & io_in2;
  assign T_194 = T_191 ? T_192 : 64'h0;
  assign logic$ = T_188 | T_194;
  assign T_195 = io_fn == 4'h2;
  assign T_196 = io_fn == 4'h3;
  assign T_197 = T_195 | T_196;
  assign T_198 = io_fn >= 4'hc;
  assign T_199 = T_197 | T_198;
  assign T_200 = T_199 & io_cmp_out;
  assign GEN_24 = {{63'd0}, T_200};
  assign T_201 = GEN_24 | logic$;
  assign shift_logic = T_201 | shout;
  assign T_202 = io_fn == 4'h0;
  assign T_203 = io_fn == 4'ha;
  assign T_204 = T_202 | T_203;
  assign out = T_204 ? io_adder_out : shift_logic;
  assign T_205 = io_dw == 1'h0;
  assign T_206 = out[31];
  assign T_210 = T_206 ? 32'hffffffff : 32'h0;
  assign T_211 = out[31:0];
  assign T_212 = {T_210,T_211};
  assign GEN_0 = T_205 ? T_212 : out;
endmodule
module MulDiv(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [3:0] io_req_bits_fn,
  input   io_req_bits_dw,
  input  [63:0] io_req_bits_in1,
  input  [63:0] io_req_bits_in2,
  input  [4:0] io_req_bits_tag,
  input   io_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [63:0] io_resp_bits_data,
  output [4:0] io_resp_bits_tag
);
  reg [2:0] state;
  reg [31:0] GEN_14;
  reg [3:0] req_fn;
  reg [31:0] GEN_15;
  reg  req_dw;
  reg [31:0] GEN_36;
  reg [63:0] req_in1;
  reg [63:0] GEN_37;
  reg [63:0] req_in2;
  reg [63:0] GEN_38;
  reg [4:0] req_tag;
  reg [31:0] GEN_39;
  reg [6:0] count;
  reg [31:0] GEN_40;
  reg  neg_out;
  reg [31:0] GEN_41;
  reg  isMul;
  reg [31:0] GEN_42;
  reg  isHi;
  reg [31:0] GEN_43;
  reg [64:0] divisor;
  reg [95:0] GEN_44;
  reg [129:0] remainder;
  reg [159:0] GEN_45;
  wire [3:0] T_62;
  wire  T_64;
  wire [3:0] T_66;
  wire  T_68;
  wire  T_71;
  wire [3:0] T_73;
  wire  T_75;
  wire [3:0] T_77;
  wire  T_79;
  wire  T_82;
  wire  T_83;
  wire [3:0] T_85;
  wire  T_87;
  wire [3:0] T_89;
  wire  T_91;
  wire  T_94;
  wire  T_95;
  wire  T_100;
  wire  T_102;
  wire  T_103;
  wire  T_104;
  wire  lhs_sign;
  wire [31:0] T_108;
  wire [31:0] T_109;
  wire [31:0] T_110;
  wire [31:0] T_111;
  wire [63:0] lhs_in;
  wire  T_115;
  wire  T_116;
  wire  T_117;
  wire  rhs_sign;
  wire [31:0] T_121;
  wire [31:0] T_122;
  wire [31:0] T_123;
  wire [31:0] T_124;
  wire [63:0] rhs_in;
  wire [64:0] T_125;
  wire [65:0] T_127;
  wire [64:0] subtractor;
  wire  less;
  wire [63:0] T_128;
  wire [64:0] T_130;
  wire [63:0] negated_remainder;
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire [129:0] GEN_0;
  wire  T_134;
  wire  T_135;
  wire [64:0] GEN_1;
  wire [129:0] GEN_2;
  wire [64:0] GEN_3;
  wire [2:0] GEN_4;
  wire  T_136;
  wire [129:0] GEN_5;
  wire [2:0] GEN_6;
  wire  T_137;
  wire [63:0] T_138;
  wire [2:0] T_139;
  wire [129:0] GEN_7;
  wire [2:0] GEN_8;
  wire  T_140;
  wire  T_141;
  wire [64:0] T_142;
  wire [128:0] T_144;
  wire [63:0] T_145;
  wire [64:0] T_146;
  wire [64:0] T_147;
  wire [64:0] T_148;
  wire  T_149;
  wire [64:0] GEN_34;
  wire [65:0] T_150;
  wire [65:0] GEN_35;
  wire [66:0] T_151;
  wire [65:0] T_152;
  wire [65:0] T_153;
  wire [62:0] T_154;
  wire [65:0] T_155;
  wire [128:0] T_156;
  wire  T_171;
  wire [64:0] T_185;
  wire [63:0] T_187;
  wire [128:0] T_188;
  wire [64:0] T_189;
  wire [63:0] T_191;
  wire [65:0] T_192;
  wire [129:0] T_193;
  wire [7:0] T_195;
  wire [6:0] T_196;
  wire  T_198;
  wire [2:0] T_200;
  wire [2:0] GEN_9;
  wire [129:0] GEN_10;
  wire [6:0] GEN_11;
  wire [2:0] GEN_12;
  wire  T_203;
  wire  T_204;
  wire  T_206;
  wire [2:0] T_208;
  wire [2:0] GEN_13;
  wire [63:0] T_212;
  wire [63:0] T_213;
  wire [63:0] T_214;
  wire  T_217;
  wire [127:0] T_218;
  wire [128:0] T_219;
  wire  T_665;
  wire  T_682;
  wire  T_685;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [6:0] GEN_18;
  wire [129:0] GEN_19;
  wire  GEN_20;
  wire  T_687;
  wire  T_688;
  wire [2:0] GEN_21;
  wire  T_689;
  wire  T_691;
  wire  T_692;
  wire  T_693;
  wire [2:0] T_694;
  wire  T_698;
  wire  T_699;
  wire  T_700;
  wire [64:0] T_701;
  wire [2:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [6:0] GEN_25;
  wire  GEN_26;
  wire [64:0] GEN_27;
  wire [129:0] GEN_28;
  wire [3:0] GEN_29;
  wire  GEN_30;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [4:0] GEN_33;
  wire  T_703;
  wire  T_705;
  wire [31:0] T_709;
  wire [31:0] T_710;
  wire [63:0] T_711;
  wire [63:0] T_713;
  wire  T_714;
  wire  T_715;
  assign io_req_ready = T_715;
  assign io_resp_valid = T_714;
  assign io_resp_bits_data = T_713;
  assign io_resp_bits_tag = req_tag;
  assign T_62 = io_req_bits_fn & 4'h4;
  assign T_64 = T_62 == 4'h0;
  assign T_66 = io_req_bits_fn & 4'h8;
  assign T_68 = T_66 == 4'h8;
  assign T_71 = T_64 | T_68;
  assign T_73 = io_req_bits_fn & 4'h5;
  assign T_75 = T_73 == 4'h1;
  assign T_77 = io_req_bits_fn & 4'h2;
  assign T_79 = T_77 == 4'h2;
  assign T_82 = T_75 | T_79;
  assign T_83 = T_82 | T_68;
  assign T_85 = io_req_bits_fn & 4'h9;
  assign T_87 = T_85 == 4'h0;
  assign T_89 = io_req_bits_fn & 4'h3;
  assign T_91 = T_89 == 4'h0;
  assign T_94 = T_87 | T_64;
  assign T_95 = T_94 | T_91;
  assign T_100 = io_req_bits_dw == 1'h0;
  assign T_102 = io_req_bits_in1[31];
  assign T_103 = io_req_bits_in1[63];
  assign T_104 = T_100 ? T_102 : T_103;
  assign lhs_sign = T_95 & T_104;
  assign T_108 = lhs_sign ? 32'hffffffff : 32'h0;
  assign T_109 = io_req_bits_in1[63:32];
  assign T_110 = T_100 ? T_108 : T_109;
  assign T_111 = io_req_bits_in1[31:0];
  assign lhs_in = {T_110,T_111};
  assign T_115 = io_req_bits_in2[31];
  assign T_116 = io_req_bits_in2[63];
  assign T_117 = T_100 ? T_115 : T_116;
  assign rhs_sign = T_94 & T_117;
  assign T_121 = rhs_sign ? 32'hffffffff : 32'h0;
  assign T_122 = io_req_bits_in2[63:32];
  assign T_123 = T_100 ? T_121 : T_122;
  assign T_124 = io_req_bits_in2[31:0];
  assign rhs_in = {T_123,T_124};
  assign T_125 = remainder[128:64];
  assign T_127 = T_125 - divisor;
  assign subtractor = T_127[64:0];
  assign less = subtractor[64];
  assign T_128 = remainder[63:0];
  assign T_130 = 64'h0 - T_128;
  assign negated_remainder = T_130[63:0];
  assign T_131 = state == 3'h1;
  assign T_132 = remainder[63];
  assign T_133 = T_132 | isMul;
  assign GEN_0 = T_133 ? {{66'd0}, negated_remainder} : remainder;
  assign T_134 = divisor[63];
  assign T_135 = T_134 | isMul;
  assign GEN_1 = T_135 ? subtractor : divisor;
  assign GEN_2 = T_131 ? GEN_0 : remainder;
  assign GEN_3 = T_131 ? GEN_1 : divisor;
  assign GEN_4 = T_131 ? 3'h2 : state;
  assign T_136 = state == 3'h4;
  assign GEN_5 = T_136 ? {{66'd0}, negated_remainder} : GEN_2;
  assign GEN_6 = T_136 ? 3'h5 : GEN_4;
  assign T_137 = state == 3'h3;
  assign T_138 = remainder[128:65];
  assign T_139 = neg_out ? 3'h4 : 3'h5;
  assign GEN_7 = T_137 ? {{66'd0}, T_138} : GEN_5;
  assign GEN_8 = T_137 ? T_139 : GEN_6;
  assign T_140 = state == 3'h2;
  assign T_141 = T_140 & isMul;
  assign T_142 = remainder[129:65];
  assign T_144 = {T_142,T_128};
  assign T_145 = T_144[63:0];
  assign T_146 = T_144[128:64];
  assign T_147 = $signed(T_146);
  assign T_148 = $signed(divisor);
  assign T_149 = T_145[0];
  assign GEN_34 = {{64'd0}, T_149};
  assign T_150 = $signed(T_148) * $signed({1'b0,GEN_34});
  assign GEN_35 = {{1{T_147[64]}},T_147};
  assign T_151 = $signed(T_150) + $signed(GEN_35);
  assign T_152 = T_151[65:0];
  assign T_153 = $signed(T_152);
  assign T_154 = T_145[63:1];
  assign T_155 = $unsigned(T_153);
  assign T_156 = {T_155,T_154};
  assign T_171 = isHi == 1'h0;
  assign T_185 = T_156[128:64];
  assign T_187 = T_156[63:0];
  assign T_188 = {T_185,T_187};
  assign T_189 = T_188[128:64];
  assign T_191 = T_188[63:0];
  assign T_192 = {T_189,1'h0};
  assign T_193 = {T_192,T_191};
  assign T_195 = count + 7'h1;
  assign T_196 = T_195[6:0];
  assign T_198 = count == 7'h3f;
  assign T_200 = isHi ? 3'h3 : 3'h5;
  assign GEN_9 = T_198 ? T_200 : GEN_8;
  assign GEN_10 = T_141 ? T_193 : GEN_7;
  assign GEN_11 = T_141 ? T_196 : count;
  assign GEN_12 = T_141 ? GEN_9 : GEN_8;
  assign T_203 = isMul == 1'h0;
  assign T_204 = T_140 & T_203;
  assign T_206 = count == 7'h40;
  assign T_208 = isHi ? 3'h3 : T_139;
  assign GEN_13 = T_206 ? T_208 : GEN_12;
  assign T_212 = remainder[127:64];
  assign T_213 = subtractor[63:0];
  assign T_214 = less ? T_212 : T_213;
  assign T_217 = less == 1'h0;
  assign T_218 = {T_214,T_128};
  assign T_219 = {T_218,T_217};
  assign T_665 = count == 7'h0;
  assign T_682 = T_665 & T_217;
  assign T_685 = T_682 & T_171;
  assign GEN_16 = T_685 ? 1'h0 : neg_out;
  assign GEN_17 = T_204 ? GEN_13 : GEN_12;
  assign GEN_18 = T_204 ? T_196 : GEN_11;
  assign GEN_19 = T_204 ? {{1'd0}, T_219} : GEN_10;
  assign GEN_20 = T_204 ? GEN_16 : neg_out;
  assign T_687 = io_resp_ready & io_resp_valid;
  assign T_688 = T_687 | io_kill;
  assign GEN_21 = T_688 ? 3'h0 : GEN_17;
  assign T_689 = io_req_ready & io_req_valid;
  assign T_691 = T_71 == 1'h0;
  assign T_692 = rhs_sign & T_691;
  assign T_693 = lhs_sign | T_692;
  assign T_694 = T_693 ? 3'h1 : 3'h2;
  assign T_698 = lhs_sign != rhs_sign;
  assign T_699 = T_83 ? lhs_sign : T_698;
  assign T_700 = T_691 & T_699;
  assign T_701 = {rhs_sign,rhs_in};
  assign GEN_22 = T_689 ? T_694 : GEN_21;
  assign GEN_23 = T_689 ? T_71 : isMul;
  assign GEN_24 = T_689 ? T_83 : isHi;
  assign GEN_25 = T_689 ? 7'h0 : GEN_18;
  assign GEN_26 = T_689 ? T_700 : GEN_20;
  assign GEN_27 = T_689 ? T_701 : GEN_3;
  assign GEN_28 = T_689 ? {{66'd0}, lhs_in} : GEN_19;
  assign GEN_29 = T_689 ? io_req_bits_fn : req_fn;
  assign GEN_30 = T_689 ? io_req_bits_dw : req_dw;
  assign GEN_31 = T_689 ? io_req_bits_in1 : req_in1;
  assign GEN_32 = T_689 ? io_req_bits_in2 : req_in2;
  assign GEN_33 = T_689 ? io_req_bits_tag : req_tag;
  assign T_703 = req_dw == 1'h0;
  assign T_705 = remainder[31];
  assign T_709 = T_705 ? 32'hffffffff : 32'h0;
  assign T_710 = remainder[31:0];
  assign T_711 = {T_709,T_710};
  assign T_713 = T_703 ? T_711 : T_128;
  assign T_714 = state == 3'h5;
  assign T_715 = state == 3'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_14 = {1{$random}};
  state = GEN_14[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_15 = {1{$random}};
  req_fn = GEN_15[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  req_dw = GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {2{$random}};
  req_in1 = GEN_37[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {2{$random}};
  req_in2 = GEN_38[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  req_tag = GEN_39[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  count = GEN_40[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  neg_out = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  isMul = GEN_42[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  isHi = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {3{$random}};
  divisor = GEN_44[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {5{$random}};
  remainder = GEN_45[129:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      if(T_689) begin
        if(T_693) begin
          state <= 3'h1;
        end else begin
          state <= 3'h2;
        end
      end else begin
        if(T_688) begin
          state <= 3'h0;
        end else begin
          if(T_204) begin
            if(T_206) begin
              if(isHi) begin
                state <= 3'h3;
              end else begin
                if(neg_out) begin
                  state <= 3'h4;
                end else begin
                  state <= 3'h5;
                end
              end
            end else begin
              if(T_141) begin
                if(T_198) begin
                  if(isHi) begin
                    state <= 3'h3;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_137) begin
                    if(neg_out) begin
                      state <= 3'h4;
                    end else begin
                      state <= 3'h5;
                    end
                  end else begin
                    if(T_136) begin
                      state <= 3'h5;
                    end else begin
                      if(T_131) begin
                        state <= 3'h2;
                      end
                    end
                  end
                end
              end else begin
                if(T_137) begin
                  if(neg_out) begin
                    state <= 3'h4;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_136) begin
                    state <= 3'h5;
                  end else begin
                    if(T_131) begin
                      state <= 3'h2;
                    end
                  end
                end
              end
            end
          end else begin
            if(T_141) begin
              if(T_198) begin
                if(isHi) begin
                  state <= 3'h3;
                end else begin
                  state <= 3'h5;
                end
              end else begin
                if(T_137) begin
                  if(neg_out) begin
                    state <= 3'h4;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_136) begin
                    state <= 3'h5;
                  end else begin
                    if(T_131) begin
                      state <= 3'h2;
                    end
                  end
                end
              end
            end else begin
              if(T_137) begin
                state <= T_139;
              end else begin
                if(T_136) begin
                  state <= 3'h5;
                end else begin
                  if(T_131) begin
                    state <= 3'h2;
                  end
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_fn <= io_req_bits_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_dw <= io_req_bits_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_in1 <= io_req_bits_in1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_in2 <= io_req_bits_in2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        count <= 7'h0;
      end else begin
        if(T_204) begin
          count <= T_196;
        end else begin
          if(T_141) begin
            count <= T_196;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        neg_out <= T_700;
      end else begin
        if(T_204) begin
          if(T_685) begin
            neg_out <= 1'h0;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        isMul <= T_71;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        isHi <= T_83;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        divisor <= T_701;
      end else begin
        if(T_131) begin
          if(T_135) begin
            divisor <= subtractor;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        remainder <= {{66'd0}, lhs_in};
      end else begin
        if(T_204) begin
          remainder <= {{1'd0}, T_219};
        end else begin
          if(T_141) begin
            remainder <= T_193;
          end else begin
            if(T_137) begin
              remainder <= {{66'd0}, T_138};
            end else begin
              if(T_136) begin
                remainder <= {{66'd0}, negated_remainder};
              end else begin
                if(T_131) begin
                  if(T_133) begin
                    remainder <= {{66'd0}, negated_remainder};
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module Rocket(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip,
  output  io_imem_req_valid,
  output [39:0] io_imem_req_bits_pc,
  output  io_imem_req_bits_speculative,
  output  io_imem_resp_ready,
  input   io_imem_resp_valid,
  input   io_imem_resp_bits_btb_valid,
  input   io_imem_resp_bits_btb_bits_taken,
  input  [1:0] io_imem_resp_bits_btb_bits_mask,
  input   io_imem_resp_bits_btb_bits_bridx,
  input  [38:0] io_imem_resp_bits_btb_bits_target,
  input   io_imem_resp_bits_btb_bits_entry,
  input   io_imem_resp_bits_btb_bits_bht_history,
  input  [1:0] io_imem_resp_bits_btb_bits_bht_value,
  input  [39:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data,
  input  [1:0] io_imem_resp_bits_mask,
  input   io_imem_resp_bits_xcpt_if,
  input   io_imem_resp_bits_replay,
  output  io_imem_btb_update_valid,
  output  io_imem_btb_update_bits_prediction_valid,
  output  io_imem_btb_update_bits_prediction_bits_taken,
  output [1:0] io_imem_btb_update_bits_prediction_bits_mask,
  output  io_imem_btb_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_btb_update_bits_prediction_bits_target,
  output  io_imem_btb_update_bits_prediction_bits_entry,
  output  io_imem_btb_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
  output [38:0] io_imem_btb_update_bits_pc,
  output [38:0] io_imem_btb_update_bits_target,
  output  io_imem_btb_update_bits_taken,
  output  io_imem_btb_update_bits_isValid,
  output  io_imem_btb_update_bits_isJump,
  output  io_imem_btb_update_bits_isReturn,
  output [38:0] io_imem_btb_update_bits_br_pc,
  output  io_imem_bht_update_valid,
  output  io_imem_bht_update_bits_prediction_valid,
  output  io_imem_bht_update_bits_prediction_bits_taken,
  output [1:0] io_imem_bht_update_bits_prediction_bits_mask,
  output  io_imem_bht_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_bht_update_bits_prediction_bits_target,
  output  io_imem_bht_update_bits_prediction_bits_entry,
  output  io_imem_bht_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
  output [38:0] io_imem_bht_update_bits_pc,
  output  io_imem_bht_update_bits_taken,
  output  io_imem_bht_update_bits_mispredict,
  output  io_imem_ras_update_valid,
  output  io_imem_ras_update_bits_isCall,
  output  io_imem_ras_update_bits_isReturn,
  output [38:0] io_imem_ras_update_bits_returnAddr,
  output  io_imem_ras_update_bits_prediction_valid,
  output  io_imem_ras_update_bits_prediction_bits_taken,
  output [1:0] io_imem_ras_update_bits_prediction_bits_mask,
  output  io_imem_ras_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_ras_update_bits_prediction_bits_target,
  output  io_imem_ras_update_bits_prediction_bits_entry,
  output  io_imem_ras_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
  output  io_imem_flush_icache,
  output  io_imem_flush_tlb,
  input  [39:0] io_imem_npc,
  input   io_dmem_req_ready,
  output  io_dmem_req_valid,
  output [39:0] io_dmem_req_bits_addr,
  output [5:0] io_dmem_req_bits_tag,
  output [4:0] io_dmem_req_bits_cmd,
  output [2:0] io_dmem_req_bits_typ,
  output  io_dmem_req_bits_phys,
  output [63:0] io_dmem_req_bits_data,
  output  io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data,
  input   io_dmem_s2_nack,
  input   io_dmem_resp_valid,
  input  [39:0] io_dmem_resp_bits_addr,
  input  [5:0] io_dmem_resp_bits_tag,
  input  [4:0] io_dmem_resp_bits_cmd,
  input  [2:0] io_dmem_resp_bits_typ,
  input  [63:0] io_dmem_resp_bits_data,
  input   io_dmem_resp_bits_replay,
  input   io_dmem_resp_bits_has_data,
  input  [63:0] io_dmem_resp_bits_data_word_bypass,
  input  [63:0] io_dmem_resp_bits_store_data,
  input   io_dmem_replay_next,
  input   io_dmem_xcpt_ma_ld,
  input   io_dmem_xcpt_ma_st,
  input   io_dmem_xcpt_pf_ld,
  input   io_dmem_xcpt_pf_st,
  output  io_dmem_invalidate_lr,
  input   io_dmem_ordered,
  output [6:0] io_ptw_ptbr_asid,
  output [37:0] io_ptw_ptbr_ppn,
  output  io_ptw_invalidate,
  output  io_ptw_status_debug,
  output [1:0] io_ptw_status_prv,
  output  io_ptw_status_sd,
  output [30:0] io_ptw_status_zero3,
  output  io_ptw_status_sd_rv32,
  output [1:0] io_ptw_status_zero2,
  output [4:0] io_ptw_status_vm,
  output [3:0] io_ptw_status_zero1,
  output  io_ptw_status_mxr,
  output  io_ptw_status_pum,
  output  io_ptw_status_mprv,
  output [1:0] io_ptw_status_xs,
  output [1:0] io_ptw_status_fs,
  output [1:0] io_ptw_status_mpp,
  output [1:0] io_ptw_status_hpp,
  output  io_ptw_status_spp,
  output  io_ptw_status_mpie,
  output  io_ptw_status_hpie,
  output  io_ptw_status_spie,
  output  io_ptw_status_upie,
  output  io_ptw_status_mie,
  output  io_ptw_status_hie,
  output  io_ptw_status_sie,
  output  io_ptw_status_uie,
  output [31:0] io_fpu_inst,
  output [63:0] io_fpu_fromint_data,
  output [2:0] io_fpu_fcsr_rm,
  input   io_fpu_fcsr_flags_valid,
  input  [4:0] io_fpu_fcsr_flags_bits,
  input  [63:0] io_fpu_store_data,
  input  [63:0] io_fpu_toint_data,
  output  io_fpu_dmem_resp_val,
  output [2:0] io_fpu_dmem_resp_type,
  output [4:0] io_fpu_dmem_resp_tag,
  output [63:0] io_fpu_dmem_resp_data,
  output  io_fpu_valid,
  input   io_fpu_fcsr_rdy,
  input   io_fpu_nack_mem,
  input   io_fpu_illegal_rm,
  output  io_fpu_killx,
  output  io_fpu_killm,
  input  [4:0] io_fpu_dec_cmd,
  input   io_fpu_dec_ldst,
  input   io_fpu_dec_wen,
  input   io_fpu_dec_ren1,
  input   io_fpu_dec_ren2,
  input   io_fpu_dec_ren3,
  input   io_fpu_dec_swap12,
  input   io_fpu_dec_swap23,
  input   io_fpu_dec_single,
  input   io_fpu_dec_fromint,
  input   io_fpu_dec_toint,
  input   io_fpu_dec_fastpipe,
  input   io_fpu_dec_fma,
  input   io_fpu_dec_div,
  input   io_fpu_dec_sqrt,
  input   io_fpu_dec_round,
  input   io_fpu_dec_wflags,
  input   io_fpu_sboard_set,
  input   io_fpu_sboard_clr,
  input  [4:0] io_fpu_sboard_clra,
  input   io_fpu_cp_req_ready,
  output  io_fpu_cp_req_valid,
  output [4:0] io_fpu_cp_req_bits_cmd,
  output  io_fpu_cp_req_bits_ldst,
  output  io_fpu_cp_req_bits_wen,
  output  io_fpu_cp_req_bits_ren1,
  output  io_fpu_cp_req_bits_ren2,
  output  io_fpu_cp_req_bits_ren3,
  output  io_fpu_cp_req_bits_swap12,
  output  io_fpu_cp_req_bits_swap23,
  output  io_fpu_cp_req_bits_single,
  output  io_fpu_cp_req_bits_fromint,
  output  io_fpu_cp_req_bits_toint,
  output  io_fpu_cp_req_bits_fastpipe,
  output  io_fpu_cp_req_bits_fma,
  output  io_fpu_cp_req_bits_div,
  output  io_fpu_cp_req_bits_sqrt,
  output  io_fpu_cp_req_bits_round,
  output  io_fpu_cp_req_bits_wflags,
  output [2:0] io_fpu_cp_req_bits_rm,
  output [1:0] io_fpu_cp_req_bits_typ,
  output [64:0] io_fpu_cp_req_bits_in1,
  output [64:0] io_fpu_cp_req_bits_in2,
  output [64:0] io_fpu_cp_req_bits_in3,
  output  io_fpu_cp_resp_ready,
  input   io_fpu_cp_resp_valid,
  input  [64:0] io_fpu_cp_resp_bits_data,
  input  [4:0] io_fpu_cp_resp_bits_exc,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [63:0] io_rocc_cmd_bits_rs1,
  output [63:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_cmd_bits_status_debug,
  output [1:0] io_rocc_cmd_bits_status_prv,
  output  io_rocc_cmd_bits_status_sd,
  output [30:0] io_rocc_cmd_bits_status_zero3,
  output  io_rocc_cmd_bits_status_sd_rv32,
  output [1:0] io_rocc_cmd_bits_status_zero2,
  output [4:0] io_rocc_cmd_bits_status_vm,
  output [3:0] io_rocc_cmd_bits_status_zero1,
  output  io_rocc_cmd_bits_status_mxr,
  output  io_rocc_cmd_bits_status_pum,
  output  io_rocc_cmd_bits_status_mprv,
  output [1:0] io_rocc_cmd_bits_status_xs,
  output [1:0] io_rocc_cmd_bits_status_fs,
  output [1:0] io_rocc_cmd_bits_status_mpp,
  output [1:0] io_rocc_cmd_bits_status_hpp,
  output  io_rocc_cmd_bits_status_spp,
  output  io_rocc_cmd_bits_status_mpie,
  output  io_rocc_cmd_bits_status_hpie,
  output  io_rocc_cmd_bits_status_spie,
  output  io_rocc_cmd_bits_status_upie,
  output  io_rocc_cmd_bits_status_mie,
  output  io_rocc_cmd_bits_status_hie,
  output  io_rocc_cmd_bits_status_sie,
  output  io_rocc_cmd_bits_status_uie,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [63:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [39:0] io_rocc_mem_req_bits_addr,
  input  [5:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [63:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [63:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [39:0] io_rocc_mem_resp_bits_addr,
  output [5:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [63:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [63:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [63:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input   io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [10:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output  io_rocc_autl_grant_bits_client_xact_id,
  output [1:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception
);
  reg  ex_ctrl_legal;
  reg [31:0] GEN_270;
  reg  ex_ctrl_fp;
  reg [31:0] GEN_271;
  reg  ex_ctrl_rocc;
  reg [31:0] GEN_272;
  reg  ex_ctrl_branch;
  reg [31:0] GEN_273;
  reg  ex_ctrl_jal;
  reg [31:0] GEN_274;
  reg  ex_ctrl_jalr;
  reg [31:0] GEN_275;
  reg  ex_ctrl_rxs2;
  reg [31:0] GEN_276;
  reg  ex_ctrl_rxs1;
  reg [31:0] GEN_277;
  reg [1:0] ex_ctrl_sel_alu2;
  reg [31:0] GEN_278;
  reg [1:0] ex_ctrl_sel_alu1;
  reg [31:0] GEN_279;
  reg [2:0] ex_ctrl_sel_imm;
  reg [31:0] GEN_280;
  reg  ex_ctrl_alu_dw;
  reg [31:0] GEN_281;
  reg [3:0] ex_ctrl_alu_fn;
  reg [31:0] GEN_282;
  reg  ex_ctrl_mem;
  reg [31:0] GEN_283;
  reg [4:0] ex_ctrl_mem_cmd;
  reg [31:0] GEN_284;
  reg [2:0] ex_ctrl_mem_type;
  reg [31:0] GEN_285;
  reg  ex_ctrl_rfs1;
  reg [31:0] GEN_286;
  reg  ex_ctrl_rfs2;
  reg [31:0] GEN_287;
  reg  ex_ctrl_rfs3;
  reg [31:0] GEN_288;
  reg  ex_ctrl_wfd;
  reg [31:0] GEN_289;
  reg  ex_ctrl_div;
  reg [31:0] GEN_290;
  reg  ex_ctrl_wxd;
  reg [31:0] GEN_291;
  reg [2:0] ex_ctrl_csr;
  reg [31:0] GEN_292;
  reg  ex_ctrl_fence_i;
  reg [31:0] GEN_293;
  reg  ex_ctrl_fence;
  reg [31:0] GEN_294;
  reg  ex_ctrl_amo;
  reg [31:0] GEN_295;
  reg  mem_ctrl_legal;
  reg [31:0] GEN_296;
  reg  mem_ctrl_fp;
  reg [31:0] GEN_297;
  reg  mem_ctrl_rocc;
  reg [31:0] GEN_298;
  reg  mem_ctrl_branch;
  reg [31:0] GEN_299;
  reg  mem_ctrl_jal;
  reg [31:0] GEN_300;
  reg  mem_ctrl_jalr;
  reg [31:0] GEN_301;
  reg  mem_ctrl_rxs2;
  reg [31:0] GEN_302;
  reg  mem_ctrl_rxs1;
  reg [31:0] GEN_303;
  reg [1:0] mem_ctrl_sel_alu2;
  reg [31:0] GEN_304;
  reg [1:0] mem_ctrl_sel_alu1;
  reg [31:0] GEN_305;
  reg [2:0] mem_ctrl_sel_imm;
  reg [31:0] GEN_306;
  reg  mem_ctrl_alu_dw;
  reg [31:0] GEN_307;
  reg [3:0] mem_ctrl_alu_fn;
  reg [31:0] GEN_308;
  reg  mem_ctrl_mem;
  reg [31:0] GEN_309;
  reg [4:0] mem_ctrl_mem_cmd;
  reg [31:0] GEN_310;
  reg [2:0] mem_ctrl_mem_type;
  reg [31:0] GEN_311;
  reg  mem_ctrl_rfs1;
  reg [31:0] GEN_312;
  reg  mem_ctrl_rfs2;
  reg [31:0] GEN_313;
  reg  mem_ctrl_rfs3;
  reg [31:0] GEN_314;
  reg  mem_ctrl_wfd;
  reg [31:0] GEN_315;
  reg  mem_ctrl_div;
  reg [31:0] GEN_316;
  reg  mem_ctrl_wxd;
  reg [31:0] GEN_317;
  reg [2:0] mem_ctrl_csr;
  reg [31:0] GEN_318;
  reg  mem_ctrl_fence_i;
  reg [31:0] GEN_319;
  reg  mem_ctrl_fence;
  reg [31:0] GEN_320;
  reg  mem_ctrl_amo;
  reg [31:0] GEN_321;
  reg  wb_ctrl_legal;
  reg [31:0] GEN_322;
  reg  wb_ctrl_fp;
  reg [31:0] GEN_323;
  reg  wb_ctrl_rocc;
  reg [31:0] GEN_324;
  reg  wb_ctrl_branch;
  reg [31:0] GEN_325;
  reg  wb_ctrl_jal;
  reg [31:0] GEN_326;
  reg  wb_ctrl_jalr;
  reg [31:0] GEN_327;
  reg  wb_ctrl_rxs2;
  reg [31:0] GEN_328;
  reg  wb_ctrl_rxs1;
  reg [31:0] GEN_329;
  reg [1:0] wb_ctrl_sel_alu2;
  reg [31:0] GEN_330;
  reg [1:0] wb_ctrl_sel_alu1;
  reg [31:0] GEN_331;
  reg [2:0] wb_ctrl_sel_imm;
  reg [31:0] GEN_332;
  reg  wb_ctrl_alu_dw;
  reg [31:0] GEN_333;
  reg [3:0] wb_ctrl_alu_fn;
  reg [31:0] GEN_334;
  reg  wb_ctrl_mem;
  reg [31:0] GEN_335;
  reg [4:0] wb_ctrl_mem_cmd;
  reg [31:0] GEN_336;
  reg [2:0] wb_ctrl_mem_type;
  reg [31:0] GEN_337;
  reg  wb_ctrl_rfs1;
  reg [31:0] GEN_338;
  reg  wb_ctrl_rfs2;
  reg [31:0] GEN_339;
  reg  wb_ctrl_rfs3;
  reg [31:0] GEN_340;
  reg  wb_ctrl_wfd;
  reg [31:0] GEN_341;
  reg  wb_ctrl_div;
  reg [31:0] GEN_342;
  reg  wb_ctrl_wxd;
  reg [31:0] GEN_343;
  reg [2:0] wb_ctrl_csr;
  reg [31:0] GEN_344;
  reg  wb_ctrl_fence_i;
  reg [31:0] GEN_345;
  reg  wb_ctrl_fence;
  reg [31:0] GEN_346;
  reg  wb_ctrl_amo;
  reg [31:0] GEN_347;
  reg  ex_reg_xcpt_interrupt;
  reg [31:0] GEN_348;
  reg  ex_reg_valid;
  reg [31:0] GEN_349;
  reg  ex_reg_rvc;
  reg [31:0] GEN_350;
  reg  ex_reg_btb_hit;
  reg [31:0] GEN_351;
  reg  ex_reg_btb_resp_taken;
  reg [31:0] GEN_352;
  reg [1:0] ex_reg_btb_resp_mask;
  reg [31:0] GEN_353;
  reg  ex_reg_btb_resp_bridx;
  reg [31:0] GEN_354;
  reg [38:0] ex_reg_btb_resp_target;
  reg [63:0] GEN_355;
  reg  ex_reg_btb_resp_entry;
  reg [31:0] GEN_356;
  reg  ex_reg_btb_resp_bht_history;
  reg [31:0] GEN_357;
  reg [1:0] ex_reg_btb_resp_bht_value;
  reg [31:0] GEN_358;
  reg  ex_reg_xcpt;
  reg [31:0] GEN_359;
  reg  ex_reg_flush_pipe;
  reg [31:0] GEN_360;
  reg  ex_reg_load_use;
  reg [31:0] GEN_361;
  reg [63:0] ex_reg_cause;
  reg [63:0] GEN_362;
  reg  ex_reg_replay;
  reg [31:0] GEN_363;
  reg [39:0] ex_reg_pc;
  reg [63:0] GEN_364;
  reg [31:0] ex_reg_inst;
  reg [31:0] GEN_365;
  reg  mem_reg_xcpt_interrupt;
  reg [31:0] GEN_366;
  reg  mem_reg_valid;
  reg [31:0] GEN_367;
  reg  mem_reg_rvc;
  reg [31:0] GEN_368;
  reg  mem_reg_btb_hit;
  reg [31:0] GEN_369;
  reg  mem_reg_btb_resp_taken;
  reg [31:0] GEN_370;
  reg [1:0] mem_reg_btb_resp_mask;
  reg [31:0] GEN_371;
  reg  mem_reg_btb_resp_bridx;
  reg [31:0] GEN_372;
  reg [38:0] mem_reg_btb_resp_target;
  reg [63:0] GEN_373;
  reg  mem_reg_btb_resp_entry;
  reg [31:0] GEN_374;
  reg  mem_reg_btb_resp_bht_history;
  reg [31:0] GEN_375;
  reg [1:0] mem_reg_btb_resp_bht_value;
  reg [31:0] GEN_376;
  reg  mem_reg_xcpt;
  reg [31:0] GEN_377;
  reg  mem_reg_replay;
  reg [31:0] GEN_378;
  reg  mem_reg_flush_pipe;
  reg [31:0] GEN_379;
  reg [63:0] mem_reg_cause;
  reg [63:0] GEN_380;
  reg  mem_reg_slow_bypass;
  reg [31:0] GEN_381;
  reg  mem_reg_load;
  reg [31:0] GEN_382;
  reg  mem_reg_store;
  reg [31:0] GEN_383;
  reg [39:0] mem_reg_pc;
  reg [63:0] GEN_384;
  reg [31:0] mem_reg_inst;
  reg [31:0] GEN_385;
  reg [63:0] mem_reg_wdata;
  reg [63:0] GEN_386;
  reg [63:0] mem_reg_rs2;
  reg [63:0] GEN_387;
  wire  take_pc_mem;
  reg  wb_reg_valid;
  reg [31:0] GEN_388;
  reg  wb_reg_xcpt;
  reg [31:0] GEN_389;
  reg  wb_reg_replay;
  reg [31:0] GEN_390;
  reg [63:0] wb_reg_cause;
  reg [63:0] GEN_391;
  reg [39:0] wb_reg_pc;
  reg [63:0] GEN_392;
  reg [31:0] wb_reg_inst;
  reg [31:0] GEN_393;
  reg [63:0] wb_reg_wdata;
  reg [63:0] GEN_394;
  reg [63:0] wb_reg_rs2;
  reg [63:0] GEN_395;
  wire  take_pc_wb;
  wire  take_pc_mem_wb;
  wire  ibuf_clk;
  wire  ibuf_reset;
  wire  ibuf_io_imem_ready;
  wire  ibuf_io_imem_valid;
  wire  ibuf_io_imem_bits_btb_valid;
  wire  ibuf_io_imem_bits_btb_bits_taken;
  wire [1:0] ibuf_io_imem_bits_btb_bits_mask;
  wire  ibuf_io_imem_bits_btb_bits_bridx;
  wire [38:0] ibuf_io_imem_bits_btb_bits_target;
  wire  ibuf_io_imem_bits_btb_bits_entry;
  wire  ibuf_io_imem_bits_btb_bits_bht_history;
  wire [1:0] ibuf_io_imem_bits_btb_bits_bht_value;
  wire [39:0] ibuf_io_imem_bits_pc;
  wire [31:0] ibuf_io_imem_bits_data;
  wire [1:0] ibuf_io_imem_bits_mask;
  wire  ibuf_io_imem_bits_xcpt_if;
  wire  ibuf_io_imem_bits_replay;
  wire  ibuf_io_kill;
  wire [39:0] ibuf_io_pc;
  wire  ibuf_io_btb_resp_taken;
  wire [1:0] ibuf_io_btb_resp_mask;
  wire  ibuf_io_btb_resp_bridx;
  wire [38:0] ibuf_io_btb_resp_target;
  wire  ibuf_io_btb_resp_entry;
  wire  ibuf_io_btb_resp_bht_history;
  wire [1:0] ibuf_io_btb_resp_bht_value;
  wire  ibuf_io_inst_0_ready;
  wire  ibuf_io_inst_0_valid;
  wire  ibuf_io_inst_0_bits_pf0;
  wire  ibuf_io_inst_0_bits_pf1;
  wire  ibuf_io_inst_0_bits_replay;
  wire  ibuf_io_inst_0_bits_btb_hit;
  wire  ibuf_io_inst_0_bits_rvc;
  wire [31:0] ibuf_io_inst_0_bits_inst_bits;
  wire [4:0] ibuf_io_inst_0_bits_inst_rd;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs3;
  wire  id_ctrl_legal;
  wire  id_ctrl_fp;
  wire  id_ctrl_rocc;
  wire  id_ctrl_branch;
  wire  id_ctrl_jal;
  wire  id_ctrl_jalr;
  wire  id_ctrl_rxs2;
  wire  id_ctrl_rxs1;
  wire [1:0] id_ctrl_sel_alu2;
  wire [1:0] id_ctrl_sel_alu1;
  wire [2:0] id_ctrl_sel_imm;
  wire  id_ctrl_alu_dw;
  wire [3:0] id_ctrl_alu_fn;
  wire  id_ctrl_mem;
  wire [4:0] id_ctrl_mem_cmd;
  wire [2:0] id_ctrl_mem_type;
  wire  id_ctrl_rfs1;
  wire  id_ctrl_rfs2;
  wire  id_ctrl_rfs3;
  wire  id_ctrl_wfd;
  wire  id_ctrl_div;
  wire  id_ctrl_wxd;
  wire [2:0] id_ctrl_csr;
  wire  id_ctrl_fence_i;
  wire  id_ctrl_fence;
  wire  id_ctrl_amo;
  wire [31:0] T_6645;
  wire  T_6647;
  wire [31:0] T_6649;
  wire  T_6651;
  wire [31:0] T_6653;
  wire  T_6655;
  wire [31:0] T_6657;
  wire  T_6659;
  wire [31:0] T_6661;
  wire  T_6663;
  wire [31:0] T_6665;
  wire  T_6667;
  wire [31:0] T_6669;
  wire  T_6671;
  wire [31:0] T_6673;
  wire  T_6675;
  wire [31:0] T_6677;
  wire  T_6679;
  wire [31:0] T_6681;
  wire  T_6683;
  wire [31:0] T_6685;
  wire  T_6687;
  wire [31:0] T_6689;
  wire  T_6691;
  wire [31:0] T_6693;
  wire  T_6695;
  wire  T_6699;
  wire [31:0] T_6701;
  wire  T_6703;
  wire  T_6707;
  wire [31:0] T_6709;
  wire  T_6711;
  wire [31:0] T_6713;
  wire  T_6715;
  wire  T_6719;
  wire [31:0] T_6721;
  wire  T_6723;
  wire [31:0] T_6725;
  wire  T_6727;
  wire [31:0] T_6729;
  wire  T_6731;
  wire  T_6733;
  wire  T_6735;
  wire  T_6737;
  wire [31:0] T_6739;
  wire  T_6741;
  wire [31:0] T_6743;
  wire  T_6745;
  wire [31:0] T_6747;
  wire  T_6749;
  wire  T_6752;
  wire  T_6753;
  wire  T_6754;
  wire  T_6755;
  wire  T_6756;
  wire  T_6757;
  wire  T_6758;
  wire  T_6759;
  wire  T_6760;
  wire  T_6761;
  wire  T_6762;
  wire  T_6763;
  wire  T_6764;
  wire  T_6765;
  wire  T_6766;
  wire  T_6767;
  wire  T_6768;
  wire  T_6769;
  wire  T_6770;
  wire  T_6771;
  wire  T_6772;
  wire  T_6773;
  wire  T_6774;
  wire  T_6775;
  wire  T_6776;
  wire  T_6777;
  wire  T_6778;
  wire [31:0] T_6782;
  wire  T_6784;
  wire [31:0] T_6788;
  wire  T_6790;
  wire [31:0] T_6794;
  wire  T_6796;
  wire [31:0] T_6800;
  wire  T_6802;
  wire [31:0] T_6804;
  wire  T_6806;
  wire [31:0] T_6808;
  wire  T_6810;
  wire  T_6813;
  wire  T_6814;
  wire [31:0] T_6816;
  wire  T_6818;
  wire [31:0] T_6820;
  wire  T_6822;
  wire [31:0] T_6824;
  wire  T_6826;
  wire [31:0] T_6828;
  wire  T_6830;
  wire  T_6833;
  wire  T_6834;
  wire  T_6835;
  wire [31:0] T_6837;
  wire  T_6839;
  wire [31:0] T_6841;
  wire  T_6843;
  wire [31:0] T_6845;
  wire  T_6847;
  wire [31:0] T_6849;
  wire  T_6851;
  wire  T_6854;
  wire  T_6855;
  wire  T_6856;
  wire  T_6857;
  wire  T_6861;
  wire [31:0] T_6863;
  wire  T_6865;
  wire  T_6868;
  wire  T_6869;
  wire  T_6870;
  wire [1:0] T_6871;
  wire [31:0] T_6873;
  wire  T_6875;
  wire  T_6878;
  wire  T_6879;
  wire  T_6880;
  wire [31:0] T_6882;
  wire  T_6884;
  wire  T_6887;
  wire [1:0] T_6888;
  wire  T_6892;
  wire  T_6896;
  wire  T_6899;
  wire  T_6903;
  wire  T_6906;
  wire  T_6910;
  wire [31:0] T_6912;
  wire  T_6914;
  wire  T_6917;
  wire  T_6918;
  wire [1:0] T_6919;
  wire [2:0] T_6920;
  wire [31:0] T_6922;
  wire  T_6924;
  wire [31:0] T_6926;
  wire  T_6928;
  wire  T_6931;
  wire [31:0] T_6933;
  wire  T_6935;
  wire [31:0] T_6937;
  wire  T_6939;
  wire [31:0] T_6941;
  wire  T_6943;
  wire  T_6946;
  wire  T_6947;
  wire [31:0] T_6949;
  wire  T_6951;
  wire [31:0] T_6953;
  wire  T_6955;
  wire  T_6959;
  wire [31:0] T_6961;
  wire  T_6963;
  wire [31:0] T_6965;
  wire  T_6967;
  wire [31:0] T_6969;
  wire  T_6971;
  wire  T_6974;
  wire  T_6975;
  wire  T_6976;
  wire  T_6977;
  wire  T_6978;
  wire [31:0] T_6980;
  wire  T_6982;
  wire [31:0] T_6984;
  wire  T_6986;
  wire [31:0] T_6988;
  wire  T_6990;
  wire [31:0] T_6992;
  wire  T_6994;
  wire  T_6997;
  wire  T_6998;
  wire  T_6999;
  wire  T_7003;
  wire [31:0] T_7005;
  wire  T_7007;
  wire  T_7010;
  wire  T_7011;
  wire  T_7012;
  wire [1:0] T_7013;
  wire [1:0] T_7014;
  wire [3:0] T_7015;
  wire [31:0] T_7017;
  wire  T_7019;
  wire [31:0] T_7021;
  wire  T_7023;
  wire  T_7027;
  wire  T_7028;
  wire  T_7029;
  wire  T_7030;
  wire  T_7031;
  wire [31:0] T_7033;
  wire  T_7035;
  wire [31:0] T_7037;
  wire  T_7039;
  wire [31:0] T_7041;
  wire  T_7043;
  wire [31:0] T_7045;
  wire  T_7047;
  wire  T_7050;
  wire  T_7051;
  wire  T_7052;
  wire [31:0] T_7054;
  wire  T_7056;
  wire [31:0] T_7058;
  wire  T_7060;
  wire  T_7063;
  wire [31:0] T_7065;
  wire  T_7067;
  wire [31:0] T_7069;
  wire  T_7071;
  wire [31:0] T_7073;
  wire  T_7075;
  wire  T_7078;
  wire  T_7079;
  wire  T_7080;
  wire [31:0] T_7082;
  wire  T_7084;
  wire [1:0] T_7088;
  wire [1:0] T_7089;
  wire [2:0] T_7090;
  wire [4:0] T_7091;
  wire [31:0] T_7093;
  wire  T_7095;
  wire [31:0] T_7099;
  wire  T_7101;
  wire [31:0] T_7105;
  wire  T_7107;
  wire [1:0] T_7110;
  wire [2:0] T_7111;
  wire [31:0] T_7117;
  wire  T_7119;
  wire  T_7125;
  wire [31:0] T_7127;
  wire  T_7129;
  wire  T_7133;
  wire [31:0] T_7135;
  wire  T_7137;
  wire  T_7141;
  wire  T_7144;
  wire  T_7145;
  wire  T_7146;
  wire  T_7147;
  wire  T_7148;
  wire  T_7149;
  wire [31:0] T_7151;
  wire  T_7153;
  wire  T_7159;
  wire [31:0] T_7163;
  wire  T_7165;
  wire [1:0] T_7168;
  wire [2:0] T_7169;
  wire [31:0] T_7171;
  wire  T_7173;
  wire  T_7179;
  wire [31:0] T_7183;
  wire  T_7185;
  wire  id_load_use;
  reg  id_reg_fence;
  reg [31:0] GEN_396;
  reg [63:0] T_7192 [0:30];
  reg [63:0] GEN_397;
  wire [63:0] T_7192_T_7201_data;
  wire [4:0] T_7192_T_7201_addr;
  wire  T_7192_T_7201_en;
  reg [63:0] GEN_398;
  wire [63:0] T_7192_T_7211_data;
  wire [4:0] T_7192_T_7211_addr;
  wire  T_7192_T_7211_en;
  reg [63:0] GEN_399;
  wire [63:0] T_7192_T_7944_data;
  wire [4:0] T_7192_T_7944_addr;
  wire  T_7192_T_7944_mask;
  wire  T_7192_T_7944_en;
  wire [63:0] id_rs_0;
  wire  T_7196;
  wire [4:0] T_7199;
  wire [4:0] T_7200;
  wire [63:0] T_7202;
  wire [63:0] id_rs_1;
  wire [4:0] T_7209;
  wire [4:0] T_7210;
  wire [63:0] T_7212;
  wire  ctrl_killd;
  wire  csr_clk;
  wire  csr_reset;
  wire  csr_io_prci_reset;
  wire  csr_io_prci_id;
  wire  csr_io_prci_interrupts_meip;
  wire  csr_io_prci_interrupts_seip;
  wire  csr_io_prci_interrupts_debug;
  wire  csr_io_prci_interrupts_mtip;
  wire  csr_io_prci_interrupts_msip;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [63:0] csr_io_rw_rdata;
  wire [63:0] csr_io_rw_wdata;
  wire  csr_io_csr_stall;
  wire  csr_io_csr_xcpt;
  wire  csr_io_eret;
  wire  csr_io_singleStep;
  wire  csr_io_status_debug;
  wire [1:0] csr_io_status_prv;
  wire  csr_io_status_sd;
  wire [30:0] csr_io_status_zero3;
  wire  csr_io_status_sd_rv32;
  wire [1:0] csr_io_status_zero2;
  wire [4:0] csr_io_status_vm;
  wire [3:0] csr_io_status_zero1;
  wire  csr_io_status_mxr;
  wire  csr_io_status_pum;
  wire  csr_io_status_mprv;
  wire [1:0] csr_io_status_xs;
  wire [1:0] csr_io_status_fs;
  wire [1:0] csr_io_status_mpp;
  wire [1:0] csr_io_status_hpp;
  wire  csr_io_status_spp;
  wire  csr_io_status_mpie;
  wire  csr_io_status_hpie;
  wire  csr_io_status_spie;
  wire  csr_io_status_upie;
  wire  csr_io_status_mie;
  wire  csr_io_status_hie;
  wire  csr_io_status_sie;
  wire  csr_io_status_uie;
  wire [6:0] csr_io_ptbr_asid;
  wire [37:0] csr_io_ptbr_ppn;
  wire [39:0] csr_io_evec;
  wire  csr_io_exception;
  wire  csr_io_retire;
  wire [63:0] csr_io_cause;
  wire [39:0] csr_io_pc;
  wire [39:0] csr_io_badaddr;
  wire  csr_io_fatc;
  wire [63:0] csr_io_time;
  wire [2:0] csr_io_fcsr_rm;
  wire  csr_io_fcsr_flags_valid;
  wire [4:0] csr_io_fcsr_flags_bits;
  wire  csr_io_rocc_cmd_ready;
  wire  csr_io_rocc_cmd_valid;
  wire [6:0] csr_io_rocc_cmd_bits_inst_funct;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs1;
  wire  csr_io_rocc_cmd_bits_inst_xd;
  wire  csr_io_rocc_cmd_bits_inst_xs1;
  wire  csr_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rd;
  wire [6:0] csr_io_rocc_cmd_bits_inst_opcode;
  wire [63:0] csr_io_rocc_cmd_bits_rs1;
  wire [63:0] csr_io_rocc_cmd_bits_rs2;
  wire  csr_io_rocc_cmd_bits_status_debug;
  wire [1:0] csr_io_rocc_cmd_bits_status_prv;
  wire  csr_io_rocc_cmd_bits_status_sd;
  wire [30:0] csr_io_rocc_cmd_bits_status_zero3;
  wire  csr_io_rocc_cmd_bits_status_sd_rv32;
  wire [1:0] csr_io_rocc_cmd_bits_status_zero2;
  wire [4:0] csr_io_rocc_cmd_bits_status_vm;
  wire [3:0] csr_io_rocc_cmd_bits_status_zero1;
  wire  csr_io_rocc_cmd_bits_status_mxr;
  wire  csr_io_rocc_cmd_bits_status_pum;
  wire  csr_io_rocc_cmd_bits_status_mprv;
  wire [1:0] csr_io_rocc_cmd_bits_status_xs;
  wire [1:0] csr_io_rocc_cmd_bits_status_fs;
  wire [1:0] csr_io_rocc_cmd_bits_status_mpp;
  wire [1:0] csr_io_rocc_cmd_bits_status_hpp;
  wire  csr_io_rocc_cmd_bits_status_spp;
  wire  csr_io_rocc_cmd_bits_status_mpie;
  wire  csr_io_rocc_cmd_bits_status_hpie;
  wire  csr_io_rocc_cmd_bits_status_spie;
  wire  csr_io_rocc_cmd_bits_status_upie;
  wire  csr_io_rocc_cmd_bits_status_mie;
  wire  csr_io_rocc_cmd_bits_status_hie;
  wire  csr_io_rocc_cmd_bits_status_sie;
  wire  csr_io_rocc_cmd_bits_status_uie;
  wire  csr_io_rocc_resp_ready;
  wire  csr_io_rocc_resp_valid;
  wire [4:0] csr_io_rocc_resp_bits_rd;
  wire [63:0] csr_io_rocc_resp_bits_data;
  wire  csr_io_rocc_mem_req_ready;
  wire  csr_io_rocc_mem_req_valid;
  wire [39:0] csr_io_rocc_mem_req_bits_addr;
  wire [5:0] csr_io_rocc_mem_req_bits_tag;
  wire [4:0] csr_io_rocc_mem_req_bits_cmd;
  wire [2:0] csr_io_rocc_mem_req_bits_typ;
  wire  csr_io_rocc_mem_req_bits_phys;
  wire [63:0] csr_io_rocc_mem_req_bits_data;
  wire  csr_io_rocc_mem_s1_kill;
  wire [63:0] csr_io_rocc_mem_s1_data;
  wire  csr_io_rocc_mem_s2_nack;
  wire  csr_io_rocc_mem_resp_valid;
  wire [39:0] csr_io_rocc_mem_resp_bits_addr;
  wire [5:0] csr_io_rocc_mem_resp_bits_tag;
  wire [4:0] csr_io_rocc_mem_resp_bits_cmd;
  wire [2:0] csr_io_rocc_mem_resp_bits_typ;
  wire [63:0] csr_io_rocc_mem_resp_bits_data;
  wire  csr_io_rocc_mem_resp_bits_replay;
  wire  csr_io_rocc_mem_resp_bits_has_data;
  wire [63:0] csr_io_rocc_mem_resp_bits_data_word_bypass;
  wire [63:0] csr_io_rocc_mem_resp_bits_store_data;
  wire  csr_io_rocc_mem_replay_next;
  wire  csr_io_rocc_mem_xcpt_ma_ld;
  wire  csr_io_rocc_mem_xcpt_ma_st;
  wire  csr_io_rocc_mem_xcpt_pf_ld;
  wire  csr_io_rocc_mem_xcpt_pf_st;
  wire  csr_io_rocc_mem_invalidate_lr;
  wire  csr_io_rocc_mem_ordered;
  wire  csr_io_rocc_busy;
  wire  csr_io_rocc_interrupt;
  wire  csr_io_rocc_autl_acquire_ready;
  wire  csr_io_rocc_autl_acquire_valid;
  wire [25:0] csr_io_rocc_autl_acquire_bits_addr_block;
  wire  csr_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] csr_io_rocc_autl_acquire_bits_addr_beat;
  wire  csr_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] csr_io_rocc_autl_acquire_bits_a_type;
  wire [10:0] csr_io_rocc_autl_acquire_bits_union;
  wire [63:0] csr_io_rocc_autl_acquire_bits_data;
  wire  csr_io_rocc_autl_grant_ready;
  wire  csr_io_rocc_autl_grant_valid;
  wire [2:0] csr_io_rocc_autl_grant_bits_addr_beat;
  wire  csr_io_rocc_autl_grant_bits_client_xact_id;
  wire [1:0] csr_io_rocc_autl_grant_bits_manager_xact_id;
  wire  csr_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] csr_io_rocc_autl_grant_bits_g_type;
  wire [63:0] csr_io_rocc_autl_grant_bits_data;
  wire  csr_io_rocc_fpu_req_ready;
  wire  csr_io_rocc_fpu_req_valid;
  wire [4:0] csr_io_rocc_fpu_req_bits_cmd;
  wire  csr_io_rocc_fpu_req_bits_ldst;
  wire  csr_io_rocc_fpu_req_bits_wen;
  wire  csr_io_rocc_fpu_req_bits_ren1;
  wire  csr_io_rocc_fpu_req_bits_ren2;
  wire  csr_io_rocc_fpu_req_bits_ren3;
  wire  csr_io_rocc_fpu_req_bits_swap12;
  wire  csr_io_rocc_fpu_req_bits_swap23;
  wire  csr_io_rocc_fpu_req_bits_single;
  wire  csr_io_rocc_fpu_req_bits_fromint;
  wire  csr_io_rocc_fpu_req_bits_toint;
  wire  csr_io_rocc_fpu_req_bits_fastpipe;
  wire  csr_io_rocc_fpu_req_bits_fma;
  wire  csr_io_rocc_fpu_req_bits_div;
  wire  csr_io_rocc_fpu_req_bits_sqrt;
  wire  csr_io_rocc_fpu_req_bits_round;
  wire  csr_io_rocc_fpu_req_bits_wflags;
  wire [2:0] csr_io_rocc_fpu_req_bits_rm;
  wire [1:0] csr_io_rocc_fpu_req_bits_typ;
  wire [64:0] csr_io_rocc_fpu_req_bits_in1;
  wire [64:0] csr_io_rocc_fpu_req_bits_in2;
  wire [64:0] csr_io_rocc_fpu_req_bits_in3;
  wire  csr_io_rocc_fpu_resp_ready;
  wire  csr_io_rocc_fpu_resp_valid;
  wire [64:0] csr_io_rocc_fpu_resp_bits_data;
  wire [4:0] csr_io_rocc_fpu_resp_bits_exc;
  wire  csr_io_rocc_exception;
  wire  csr_io_interrupt;
  wire [63:0] csr_io_interrupt_cause;
  wire [3:0] csr_io_bp_0_control_ttype;
  wire  csr_io_bp_0_control_dmode;
  wire [5:0] csr_io_bp_0_control_maskmax;
  wire [39:0] csr_io_bp_0_control_reserved;
  wire  csr_io_bp_0_control_action;
  wire  csr_io_bp_0_control_chain;
  wire [1:0] csr_io_bp_0_control_zero;
  wire [1:0] csr_io_bp_0_control_tmatch;
  wire  csr_io_bp_0_control_m;
  wire  csr_io_bp_0_control_h;
  wire  csr_io_bp_0_control_s;
  wire  csr_io_bp_0_control_u;
  wire  csr_io_bp_0_control_x;
  wire  csr_io_bp_0_control_w;
  wire  csr_io_bp_0_control_r;
  wire [38:0] csr_io_bp_0_address;
  wire  id_csr_en;
  wire  id_system_insn;
  wire  T_7214;
  wire  T_7215;
  wire  T_7216;
  wire  id_csr_ren;
  wire [2:0] id_csr;
  wire [11:0] id_csr_addr;
  wire  T_7220;
  wire  T_7221;
  wire [11:0] T_7351;
  wire  T_7353;
  wire [11:0] T_7355;
  wire  T_7357;
  wire  T_7360;
  wire  T_7363;
  wire  T_7364;
  wire  id_csr_flush;
  wire  T_7366;
  wire  T_7368;
  wire  T_7370;
  wire  T_7371;
  wire  T_7372;
  wire  T_7374;
  wire  T_7376;
  wire  T_7377;
  wire  id_illegal_insn;
  wire  id_amo_aq;
  wire  id_amo_rl;
  wire  T_7378;
  wire  id_fence_next;
  wire  T_7380;
  wire  id_mem_busy;
  wire  T_7386;
  wire  T_7388;
  wire  T_7389;
  wire  T_7391;
  wire  T_7392;
  wire  T_7393;
  wire  T_7394;
  wire  T_7395;
  wire  T_7396;
  wire  T_7397;
  wire  bpu_clk;
  wire  bpu_reset;
  wire  bpu_io_status_debug;
  wire [1:0] bpu_io_status_prv;
  wire  bpu_io_status_sd;
  wire [30:0] bpu_io_status_zero3;
  wire  bpu_io_status_sd_rv32;
  wire [1:0] bpu_io_status_zero2;
  wire [4:0] bpu_io_status_vm;
  wire [3:0] bpu_io_status_zero1;
  wire  bpu_io_status_mxr;
  wire  bpu_io_status_pum;
  wire  bpu_io_status_mprv;
  wire [1:0] bpu_io_status_xs;
  wire [1:0] bpu_io_status_fs;
  wire [1:0] bpu_io_status_mpp;
  wire [1:0] bpu_io_status_hpp;
  wire  bpu_io_status_spp;
  wire  bpu_io_status_mpie;
  wire  bpu_io_status_hpie;
  wire  bpu_io_status_spie;
  wire  bpu_io_status_upie;
  wire  bpu_io_status_mie;
  wire  bpu_io_status_hie;
  wire  bpu_io_status_sie;
  wire  bpu_io_status_uie;
  wire [3:0] bpu_io_bp_0_control_ttype;
  wire  bpu_io_bp_0_control_dmode;
  wire [5:0] bpu_io_bp_0_control_maskmax;
  wire [39:0] bpu_io_bp_0_control_reserved;
  wire  bpu_io_bp_0_control_action;
  wire  bpu_io_bp_0_control_chain;
  wire [1:0] bpu_io_bp_0_control_zero;
  wire [1:0] bpu_io_bp_0_control_tmatch;
  wire  bpu_io_bp_0_control_m;
  wire  bpu_io_bp_0_control_h;
  wire  bpu_io_bp_0_control_s;
  wire  bpu_io_bp_0_control_u;
  wire  bpu_io_bp_0_control_x;
  wire  bpu_io_bp_0_control_w;
  wire  bpu_io_bp_0_control_r;
  wire [38:0] bpu_io_bp_0_address;
  wire [38:0] bpu_io_pc;
  wire [38:0] bpu_io_ea;
  wire  bpu_io_xcpt_if;
  wire  bpu_io_xcpt_ld;
  wire  bpu_io_xcpt_st;
  wire  bpu_io_debug_if;
  wire  bpu_io_debug_ld;
  wire  bpu_io_debug_st;
  wire  id_xcpt_if;
  wire  T_7402;
  wire  T_7403;
  wire  T_7404;
  wire  id_xcpt;
  wire [1:0] T_7405;
  wire [1:0] T_7406;
  wire [3:0] T_7407;
  wire [63:0] id_cause;
  wire [4:0] ex_waddr;
  wire [4:0] mem_waddr;
  wire [4:0] wb_waddr;
  wire  T_7411;
  wire  T_7412;
  wire  T_7414;
  wire  T_7415;
  wire  T_7417;
  wire  T_7418;
  wire  id_bypass_src_0_1;
  wire  T_7419;
  wire  id_bypass_src_0_2;
  wire  id_bypass_src_0_3;
  wire  T_7421;
  wire  T_7422;
  wire  id_bypass_src_1_1;
  wire  T_7423;
  wire  id_bypass_src_1_2;
  wire  id_bypass_src_1_3;
  wire [63:0] bypass_mux_0;
  wire [63:0] bypass_mux_1;
  wire [63:0] bypass_mux_2;
  wire [63:0] bypass_mux_3;
  reg  ex_reg_rs_bypass_0;
  reg [31:0] GEN_400;
  reg  ex_reg_rs_bypass_1;
  reg [31:0] GEN_401;
  reg [1:0] ex_reg_rs_lsb_0;
  reg [31:0] GEN_402;
  reg [1:0] ex_reg_rs_lsb_1;
  reg [31:0] GEN_403;
  reg [61:0] ex_reg_rs_msb_0;
  reg [63:0] GEN_404;
  reg [61:0] ex_reg_rs_msb_1;
  reg [63:0] GEN_405;
  wire [63:0] T_7452;
  wire [63:0] GEN_0;
  wire [63:0] GEN_2;
  wire [63:0] GEN_3;
  wire [63:0] GEN_4;
  wire [63:0] ex_rs_0;
  wire [63:0] T_7453;
  wire [63:0] GEN_1;
  wire [63:0] GEN_5;
  wire [63:0] GEN_6;
  wire [63:0] GEN_7;
  wire [63:0] ex_rs_1;
  wire  T_7454;
  wire  T_7456;
  wire  T_7457;
  wire  T_7458;
  wire  T_7459;
  wire [10:0] T_7460;
  wire [10:0] T_7461;
  wire [10:0] T_7462;
  wire  T_7463;
  wire  T_7464;
  wire  T_7465;
  wire [7:0] T_7466;
  wire [7:0] T_7467;
  wire [7:0] T_7468;
  wire  T_7471;
  wire  T_7473;
  wire  T_7474;
  wire  T_7475;
  wire  T_7476;
  wire  T_7477;
  wire  T_7478;
  wire  T_7479;
  wire  T_7480;
  wire  T_7481;
  wire [5:0] T_7486;
  wire [5:0] T_7487;
  wire  T_7490;
  wire  T_7492;
  wire [3:0] T_7493;
  wire [3:0] T_7495;
  wire [3:0] T_7496;
  wire [3:0] T_7497;
  wire [3:0] T_7498;
  wire [3:0] T_7499;
  wire  T_7502;
  wire  T_7505;
  wire  T_7508;
  wire  T_7510;
  wire  T_7512;
  wire [9:0] T_7513;
  wire [10:0] T_7514;
  wire  T_7515;
  wire [7:0] T_7516;
  wire [8:0] T_7517;
  wire [10:0] T_7518;
  wire  T_7519;
  wire [11:0] T_7520;
  wire [20:0] T_7521;
  wire [31:0] T_7522;
  wire [31:0] ex_imm;
  wire [63:0] T_7524;
  wire [39:0] T_7525;
  wire  T_7526;
  wire [39:0] T_7527;
  wire  T_7528;
  wire [63:0] ex_op1;
  wire [63:0] T_7530;
  wire [3:0] T_7533;
  wire  T_7534;
  wire [3:0] T_7535;
  wire  T_7536;
  wire [31:0] T_7537;
  wire  T_7538;
  wire [63:0] ex_op2;
  wire  alu_clk;
  wire  alu_reset;
  wire  alu_io_dw;
  wire [3:0] alu_io_fn;
  wire [63:0] alu_io_in2;
  wire [63:0] alu_io_in1;
  wire [63:0] alu_io_out;
  wire [63:0] alu_io_adder_out;
  wire  alu_io_cmp_out;
  wire [63:0] T_7539;
  wire [63:0] T_7540;
  wire  div_clk;
  wire  div_reset;
  wire  div_io_req_ready;
  wire  div_io_req_valid;
  wire [3:0] div_io_req_bits_fn;
  wire  div_io_req_bits_dw;
  wire [63:0] div_io_req_bits_in1;
  wire [63:0] div_io_req_bits_in2;
  wire [4:0] div_io_req_bits_tag;
  wire  div_io_kill;
  wire  div_io_resp_ready;
  wire  div_io_resp_valid;
  wire [63:0] div_io_resp_bits_data;
  wire [4:0] div_io_resp_bits_tag;
  wire  T_7541;
  wire  T_7543;
  wire  T_7545;
  wire  T_7546;
  wire  T_7547;
  wire  T_7550;
  wire  T_7554;
  wire [63:0] GEN_8;
  wire  GEN_9;
  wire [1:0] GEN_10;
  wire  GEN_11;
  wire [38:0] GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [1:0] GEN_15;
  wire  T_7558;
  wire  T_7560;
  wire  T_7561;
  wire  T_7562;
  wire [1:0] GEN_16;
  wire  GEN_17;
  wire [3:0] GEN_18;
  wire  GEN_19;
  wire [1:0] GEN_20;
  wire [1:0] GEN_21;
  wire  GEN_22;
  wire  T_7564;
  wire  T_7565;
  wire  T_7566;
  wire  GEN_23;
  wire  GEN_24;
  wire  T_7569;
  wire  T_7570;
  wire  T_7571;
  wire [1:0] T_7576;
  wire [1:0] T_7577;
  wire [1:0] T_7578;
  wire  T_7580;
  wire  T_7581;
  wire [1:0] T_7582;
  wire [61:0] T_7583;
  wire [1:0] GEN_25;
  wire [61:0] GEN_26;
  wire  T_7584;
  wire  T_7585;
  wire  T_7586;
  wire [1:0] T_7591;
  wire [1:0] T_7592;
  wire [1:0] T_7593;
  wire  T_7595;
  wire  T_7596;
  wire [1:0] T_7597;
  wire [61:0] T_7598;
  wire [1:0] GEN_27;
  wire [61:0] GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire [1:0] GEN_37;
  wire [1:0] GEN_38;
  wire [2:0] GEN_39;
  wire  GEN_40;
  wire [3:0] GEN_41;
  wire  GEN_42;
  wire [4:0] GEN_43;
  wire [2:0] GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire [2:0] GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire [1:0] GEN_59;
  wire [61:0] GEN_60;
  wire  GEN_61;
  wire [1:0] GEN_62;
  wire [61:0] GEN_63;
  wire  T_7601;
  wire  T_7602;
  wire [31:0] GEN_64;
  wire [39:0] GEN_65;
  wire  T_7603;
  wire  ex_pc_valid;
  wire  T_7605;
  wire  wb_dcache_miss;
  wire  T_7607;
  wire  T_7608;
  wire  T_7610;
  wire  T_7611;
  wire  replay_ex_structural;
  wire  replay_ex_load_use;
  wire  T_7612;
  wire  T_7613;
  wire  replay_ex;
  wire  T_7614;
  wire  T_7616;
  wire  ctrl_killx;
  wire  T_7617;
  wire [2:0] T_7623_0;
  wire [2:0] T_7623_1;
  wire [2:0] T_7623_2;
  wire [2:0] T_7623_3;
  wire  T_7625;
  wire  T_7626;
  wire  T_7627;
  wire  T_7628;
  wire  T_7631;
  wire  T_7632;
  wire  T_7633;
  wire  ex_slow_bypass;
  wire  T_7634;
  wire  T_7635;
  wire  ex_xcpt;
  wire [63:0] ex_cause;
  wire  mem_br_taken;
  wire [39:0] T_7637;
  wire  T_7638;
  wire  T_7641;
  wire  T_7642;
  wire [10:0] T_7647;
  wire [7:0] T_7651;
  wire [7:0] T_7652;
  wire [7:0] T_7653;
  wire  T_7659;
  wire  T_7660;
  wire  T_7662;
  wire  T_7663;
  wire [5:0] T_7671;
  wire [3:0] T_7678;
  wire [3:0] T_7681;
  wire [9:0] T_7698;
  wire [10:0] T_7699;
  wire  T_7700;
  wire [7:0] T_7701;
  wire [8:0] T_7702;
  wire [10:0] T_7703;
  wire  T_7704;
  wire [11:0] T_7705;
  wire [20:0] T_7706;
  wire [31:0] T_7707;
  wire [31:0] T_7708;
  wire [9:0] T_7768;
  wire [10:0] T_7769;
  wire  T_7770;
  wire [7:0] T_7771;
  wire [8:0] T_7772;
  wire [20:0] T_7776;
  wire [31:0] T_7777;
  wire [31:0] T_7778;
  wire [3:0] T_7781;
  wire [31:0] T_7782;
  wire [31:0] T_7783;
  wire [39:0] GEN_171;
  wire [40:0] T_7784;
  wire [39:0] T_7785;
  wire [39:0] mem_br_target;
  wire [25:0] T_7786;
  wire [1:0] T_7787;
  wire [1:0] T_7788;
  wire  T_7790;
  wire  T_7792;
  wire  T_7793;
  wire  T_7795;
  wire [25:0] T_7796;
  wire  T_7798;
  wire  T_7801;
  wire  T_7802;
  wire  T_7804;
  wire  T_7805;
  wire  T_7806;
  wire  T_7807;
  wire [38:0] T_7808;
  wire [39:0] T_7809;
  wire [39:0] T_7810;
  wire [39:0] T_7811;
  wire [39:0] T_7813;
  wire [39:0] T_7814;
  wire [39:0] mem_npc;
  wire  T_7815;
  wire  T_7816;
  wire  T_7818;
  wire  mem_wrong_npc;
  wire  T_7820;
  wire  T_7822;
  wire [63:0] T_7823;
  wire [63:0] T_7824;
  wire [63:0] mem_int_wdata;
  wire  T_7825;
  wire  mem_cfi;
  wire  T_7827;
  wire  mem_misprediction;
  wire  T_7828;
  wire  T_7829;
  wire  T_7831;
  wire  T_7834;
  wire  T_7837;
  wire  T_7840;
  wire [63:0] GEN_66;
  wire  T_7841;
  wire  T_7842;
  wire  T_7843;
  wire  T_7845;
  wire  T_7846;
  wire  T_7847;
  wire  T_7848;
  wire  T_7849;
  wire  T_7850;
  wire  T_7851;
  wire  T_7853;
  wire  T_7857;
  wire  T_7858;
  wire  GEN_67;
  wire [1:0] GEN_68;
  wire  GEN_69;
  wire [38:0] GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire [1:0] GEN_73;
  wire  T_7859;
  wire  T_7860;
  wire [63:0] GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire [1:0] GEN_83;
  wire [1:0] GEN_84;
  wire [2:0] GEN_85;
  wire  GEN_86;
  wire [3:0] GEN_87;
  wire  GEN_88;
  wire [4:0] GEN_89;
  wire [2:0] GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire [2:0] GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire [1:0] GEN_106;
  wire  GEN_107;
  wire [38:0] GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire [1:0] GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire [31:0] GEN_114;
  wire [39:0] GEN_115;
  wire [63:0] GEN_116;
  wire [63:0] GEN_117;
  wire  T_7861;
  wire  T_7862;
  wire  mem_breakpoint;
  wire  T_7863;
  wire  T_7864;
  wire  mem_debug_breakpoint;
  wire  T_7868;
  wire  T_7870;
  wire  T_7872;
  wire  T_7874;
  wire  T_7876;
  wire  T_7878;
  wire  T_7879;
  wire  T_7880;
  wire  mem_new_xcpt;
  wire [2:0] T_7881;
  wire [2:0] T_7882;
  wire [2:0] T_7883;
  wire [2:0] T_7885;
  wire [3:0] mem_new_cause;
  wire  T_7886;
  wire  T_7887;
  wire  mem_xcpt;
  wire [63:0] mem_cause;
  wire  dcache_kill_mem;
  wire  T_7889;
  wire  fpu_kill_mem;
  wire  T_7890;
  wire  replay_mem;
  wire  T_7891;
  wire  T_7892;
  wire  T_7894;
  wire  killm_common;
  wire  T_7895;
  reg  T_7896;
  reg [31:0] GEN_406;
  wire  T_7897;
  wire  T_7898;
  wire  ctrl_killm;
  wire  T_7900;
  wire  T_7902;
  wire  T_7903;
  wire  T_7906;
  wire [63:0] GEN_118;
  wire  T_7907;
  wire  T_7908;
  wire  T_7911;
  wire  T_7912;
  wire [63:0] T_7913;
  wire [63:0] GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire [1:0] GEN_128;
  wire [1:0] GEN_129;
  wire [2:0] GEN_130;
  wire  GEN_131;
  wire [3:0] GEN_132;
  wire  GEN_133;
  wire [4:0] GEN_134;
  wire [2:0] GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire [2:0] GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire [63:0] GEN_146;
  wire [63:0] GEN_147;
  wire [31:0] GEN_148;
  wire [39:0] GEN_149;
  wire  T_7914;
  wire  wb_set_sboard;
  wire  replay_wb_common;
  wire  T_7917;
  wire  replay_wb_rocc;
  wire  replay_wb;
  wire  wb_xcpt;
  wire  T_7918;
  wire  T_7919;
  wire  T_7920;
  wire  dmem_resp_xpu;
  wire [4:0] dmem_resp_waddr;
  wire  dmem_resp_valid;
  wire  dmem_resp_replay;
  wire  T_7924;
  wire  T_7926;
  wire [63:0] ll_wdata;
  wire [4:0] ll_waddr;
  wire  T_7927;
  wire  ll_wen;
  wire  T_7928;
  wire  GEN_150;
  wire [4:0] GEN_151;
  wire  GEN_152;
  wire  T_7932;
  wire  T_7933;
  wire  T_7935;
  wire  wb_valid;
  wire  wb_wen;
  wire  rf_wen;
  wire [4:0] rf_waddr;
  wire  T_7936;
  wire  T_7937;
  wire [63:0] T_7938;
  wire [63:0] T_7939;
  wire [63:0] rf_wdata;
  wire  T_7941;
  wire [4:0] T_7943;
  wire  T_7945;
  wire [63:0] GEN_153;
  wire  T_7946;
  wire [63:0] GEN_154;
  wire [63:0] GEN_160;
  wire [63:0] GEN_161;
  wire  GEN_164;
  wire [63:0] GEN_167;
  wire [63:0] GEN_168;
  wire [25:0] T_7947;
  wire [1:0] T_7948;
  wire [1:0] T_7949;
  wire  T_7951;
  wire  T_7953;
  wire  T_7954;
  wire  T_7956;
  wire [25:0] T_7957;
  wire  T_7959;
  wire  T_7962;
  wire  T_7963;
  wire  T_7965;
  wire  T_7966;
  wire  T_7967;
  wire  T_7968;
  wire [38:0] T_7969;
  wire [39:0] T_7970;
  wire [11:0] T_7971;
  wire [2:0] T_7972;
  wire  T_7974;
  wire  T_7975;
  wire  T_7977;
  wire  T_7978;
  wire  T_7980;
  wire  T_7981;
  reg [31:0] T_7983;
  reg [31:0] GEN_407;
  wire [30:0] T_7984;
  wire [31:0] GEN_172;
  wire [31:0] T_7985;
  wire [31:0] T_7988;
  wire [31:0] T_7990;
  wire [31:0] T_7991;
  wire [31:0] T_7992;
  wire [31:0] GEN_169;
  wire [31:0] T_7994;
  wire  T_7995;
  wire  T_7996;
  wire [31:0] T_7997;
  wire  T_7998;
  wire  T_7999;
  wire [31:0] T_8000;
  wire  T_8001;
  wire  T_8002;
  wire  T_8003;
  wire  id_sboard_hazard;
  wire  T_8004;
  wire [31:0] T_8006;
  wire [31:0] T_8008;
  wire [31:0] T_8009;
  wire  T_8010;
  wire [31:0] GEN_170;
  wire  T_8011;
  wire  T_8012;
  wire  T_8013;
  wire  T_8014;
  wire  T_8015;
  wire  ex_cannot_bypass;
  wire  T_8016;
  wire  T_8017;
  wire  T_8018;
  wire  T_8019;
  wire  T_8020;
  wire  T_8021;
  wire  T_8022;
  wire  T_8023;
  wire  data_hazard_ex;
  wire  T_8025;
  wire  T_8027;
  wire  T_8028;
  wire  T_8029;
  wire  T_8031;
  wire  T_8032;
  wire  T_8033;
  wire  T_8034;
  wire  fp_data_hazard_ex;
  wire  T_8035;
  wire  T_8036;
  wire  id_ex_hazard;
  wire  T_8038;
  wire  T_8039;
  wire  T_8040;
  wire  T_8041;
  wire  T_8042;
  wire  mem_cannot_bypass;
  wire  T_8043;
  wire  T_8044;
  wire  T_8045;
  wire  T_8046;
  wire  T_8047;
  wire  T_8048;
  wire  T_8049;
  wire  T_8050;
  wire  data_hazard_mem;
  wire  T_8052;
  wire  T_8054;
  wire  T_8055;
  wire  T_8056;
  wire  T_8058;
  wire  T_8059;
  wire  T_8060;
  wire  T_8061;
  wire  fp_data_hazard_mem;
  wire  T_8062;
  wire  T_8063;
  wire  id_mem_hazard;
  wire  T_8064;
  wire  T_8065;
  wire  T_8066;
  wire  T_8067;
  wire  T_8068;
  wire  T_8069;
  wire  T_8070;
  wire  T_8071;
  wire  T_8072;
  wire  T_8073;
  wire  data_hazard_wb;
  wire  T_8075;
  wire  T_8077;
  wire  T_8078;
  wire  T_8079;
  wire  T_8081;
  wire  T_8082;
  wire  T_8083;
  wire  T_8084;
  wire  fp_data_hazard_wb;
  wire  T_8085;
  wire  T_8086;
  wire  id_wb_hazard;
  reg  dcache_blocked;
  reg [31:0] GEN_408;
  wire  T_8090;
  wire  T_8091;
  reg  rocc_blocked;
  reg [31:0] GEN_409;
  wire  T_8094;
  wire  T_8097;
  wire  T_8098;
  wire  T_8099;
  wire  T_8100;
  wire  T_8101;
  wire  T_8102;
  wire  T_8105;
  wire  T_8106;
  wire  T_8107;
  wire  T_8108;
  wire  T_8109;
  wire  ctrl_stalld;
  wire  T_8111;
  wire  T_8112;
  wire  T_8113;
  wire  T_8114;
  wire  T_8115;
  wire  T_8118;
  wire [39:0] T_8119;
  wire [39:0] T_8120;
  wire  T_8121;
  wire  T_8123;
  wire  T_8124;
  wire  T_8126;
  wire  T_8127;
  wire  T_8128;
  wire  T_8131;
  wire  T_8133;
  wire  T_8134;
  wire  T_8135;
  wire  T_8136;
  wire  T_8137;
  wire  T_8139;
  wire  T_8140;
  wire  T_8141;
  wire [4:0] T_8142;
  wire [4:0] T_8145;
  wire  T_8146;
  wire  T_8147;
  wire [1:0] T_8150;
  wire [39:0] GEN_173;
  wire [40:0] T_8151;
  wire [39:0] T_8152;
  wire [38:0] T_8153;
  wire [38:0] T_8155;
  wire [38:0] T_8156;
  wire  T_8160;
  wire  T_8164;
  wire  T_8165;
  wire  T_8168;
  wire  T_8169;
  wire  T_8170;
  wire [5:0] ex_dcache_tag;
  wire [25:0] T_8172;
  wire [1:0] T_8173;
  wire [1:0] T_8174;
  wire  T_8176;
  wire  T_8178;
  wire  T_8179;
  wire  T_8181;
  wire [25:0] T_8182;
  wire  T_8184;
  wire  T_8187;
  wire  T_8188;
  wire  T_8190;
  wire  T_8191;
  wire  T_8192;
  wire  T_8193;
  wire [38:0] T_8194;
  wire [39:0] T_8195;
  wire [63:0] T_8196;
  wire  T_8197;
  wire  T_8199;
  wire  T_8200;
  wire [1:0] T_8201;
  wire [1:0] T_8202;
  wire [3:0] T_8203;
  wire  T_8205;
  wire  T_8206;
  wire  T_8208;
  wire  T_8211;
  wire  T_8212;
  wire  T_8215;
  wire [6:0] T_8234_funct;
  wire [4:0] T_8234_rs2;
  wire [4:0] T_8234_rs1;
  wire  T_8234_xd;
  wire  T_8234_xs1;
  wire  T_8234_xs2;
  wire [4:0] T_8234_rd;
  wire [6:0] T_8234_opcode;
  wire [31:0] T_8244;
  wire [6:0] T_8245;
  wire [4:0] T_8246;
  wire  T_8247;
  wire  T_8248;
  wire  T_8249;
  wire [4:0] T_8250;
  wire [4:0] T_8251;
  wire [6:0] T_8252;
  wire [31:0] T_8253;
  wire [4:0] T_8255;
  wire [4:0] T_8256;
  reg [63:0] T_8257;
  reg [63:0] GEN_410;
  reg [63:0] T_8258;
  reg [63:0] GEN_411;
  wire [4:0] T_8259;
  reg [63:0] T_8260;
  reg [63:0] GEN_412;
  reg [63:0] T_8261;
  reg [63:0] GEN_413;
  wire  T_8263;
  wire  GEN_155;
  reg [31:0] GEN_414;
  wire [63:0] GEN_156;
  reg [63:0] GEN_415;
  wire  GEN_157;
  reg [31:0] GEN_416;
  wire [4:0] GEN_158;
  reg [31:0] GEN_417;
  wire  GEN_159;
  reg [31:0] GEN_418;
  wire  GEN_162;
  reg [31:0] GEN_419;
  wire  GEN_163;
  reg [31:0] GEN_420;
  wire  GEN_165;
  reg [31:0] GEN_421;
  wire  GEN_166;
  reg [31:0] GEN_422;
  wire  GEN_174;
  reg [31:0] GEN_423;
  wire  GEN_175;
  reg [31:0] GEN_424;
  wire  GEN_176;
  reg [31:0] GEN_425;
  wire  GEN_177;
  reg [31:0] GEN_426;
  wire  GEN_178;
  reg [31:0] GEN_427;
  wire  GEN_179;
  reg [31:0] GEN_428;
  wire  GEN_180;
  reg [31:0] GEN_429;
  wire  GEN_181;
  reg [31:0] GEN_430;
  wire  GEN_182;
  reg [31:0] GEN_431;
  wire  GEN_183;
  reg [31:0] GEN_432;
  wire  GEN_184;
  reg [31:0] GEN_433;
  wire [2:0] GEN_185;
  reg [31:0] GEN_434;
  wire [1:0] GEN_186;
  reg [31:0] GEN_435;
  wire [64:0] GEN_187;
  reg [95:0] GEN_436;
  wire [64:0] GEN_188;
  reg [95:0] GEN_437;
  wire [64:0] GEN_189;
  reg [95:0] GEN_438;
  wire  GEN_190;
  reg [31:0] GEN_439;
  wire  GEN_191;
  reg [31:0] GEN_440;
  wire  GEN_192;
  reg [31:0] GEN_441;
  wire  GEN_193;
  reg [31:0] GEN_442;
  wire  GEN_194;
  reg [31:0] GEN_443;
  wire [39:0] GEN_195;
  reg [63:0] GEN_444;
  wire [5:0] GEN_196;
  reg [31:0] GEN_445;
  wire [4:0] GEN_197;
  reg [31:0] GEN_446;
  wire [2:0] GEN_198;
  reg [31:0] GEN_447;
  wire [63:0] GEN_199;
  reg [63:0] GEN_448;
  wire  GEN_200;
  reg [31:0] GEN_449;
  wire  GEN_201;
  reg [31:0] GEN_450;
  wire [63:0] GEN_202;
  reg [63:0] GEN_451;
  wire [63:0] GEN_203;
  reg [63:0] GEN_452;
  wire  GEN_204;
  reg [31:0] GEN_453;
  wire  GEN_205;
  reg [31:0] GEN_454;
  wire  GEN_206;
  reg [31:0] GEN_455;
  wire  GEN_207;
  reg [31:0] GEN_456;
  wire  GEN_208;
  reg [31:0] GEN_457;
  wire  GEN_209;
  reg [31:0] GEN_458;
  wire  GEN_210;
  reg [31:0] GEN_459;
  wire  GEN_211;
  reg [31:0] GEN_460;
  wire [2:0] GEN_212;
  reg [31:0] GEN_461;
  wire  GEN_213;
  reg [31:0] GEN_462;
  wire [1:0] GEN_214;
  reg [31:0] GEN_463;
  wire  GEN_215;
  reg [31:0] GEN_464;
  wire [3:0] GEN_216;
  reg [31:0] GEN_465;
  wire [63:0] GEN_217;
  reg [63:0] GEN_466;
  wire  GEN_218;
  reg [31:0] GEN_467;
  wire  GEN_219;
  reg [31:0] GEN_468;
  wire [64:0] GEN_220;
  reg [95:0] GEN_469;
  wire [4:0] GEN_221;
  reg [31:0] GEN_470;
  wire  GEN_222;
  reg [31:0] GEN_471;
  wire  GEN_223;
  reg [31:0] GEN_472;
  wire [4:0] GEN_224;
  reg [31:0] GEN_473;
  wire [63:0] GEN_225;
  reg [63:0] GEN_474;
  wire  GEN_226;
  reg [31:0] GEN_475;
  wire [39:0] GEN_227;
  reg [63:0] GEN_476;
  wire [5:0] GEN_228;
  reg [31:0] GEN_477;
  wire [4:0] GEN_229;
  reg [31:0] GEN_478;
  wire [2:0] GEN_230;
  reg [31:0] GEN_479;
  wire  GEN_231;
  reg [31:0] GEN_480;
  wire [63:0] GEN_232;
  reg [63:0] GEN_481;
  wire  GEN_233;
  reg [31:0] GEN_482;
  wire [63:0] GEN_234;
  reg [63:0] GEN_483;
  wire  GEN_235;
  reg [31:0] GEN_484;
  wire  GEN_236;
  reg [31:0] GEN_485;
  wire  GEN_237;
  reg [31:0] GEN_486;
  wire [25:0] GEN_238;
  reg [31:0] GEN_487;
  wire  GEN_239;
  reg [31:0] GEN_488;
  wire [2:0] GEN_240;
  reg [31:0] GEN_489;
  wire  GEN_241;
  reg [31:0] GEN_490;
  wire [2:0] GEN_242;
  reg [31:0] GEN_491;
  wire [10:0] GEN_243;
  reg [31:0] GEN_492;
  wire [63:0] GEN_244;
  reg [63:0] GEN_493;
  wire  GEN_245;
  reg [31:0] GEN_494;
  wire  GEN_246;
  reg [31:0] GEN_495;
  wire [4:0] GEN_247;
  reg [31:0] GEN_496;
  wire  GEN_248;
  reg [31:0] GEN_497;
  wire  GEN_249;
  reg [31:0] GEN_498;
  wire  GEN_250;
  reg [31:0] GEN_499;
  wire  GEN_251;
  reg [31:0] GEN_500;
  wire  GEN_252;
  reg [31:0] GEN_501;
  wire  GEN_253;
  reg [31:0] GEN_502;
  wire  GEN_254;
  reg [31:0] GEN_503;
  wire  GEN_255;
  reg [31:0] GEN_504;
  wire  GEN_256;
  reg [31:0] GEN_505;
  wire  GEN_257;
  reg [31:0] GEN_506;
  wire  GEN_258;
  reg [31:0] GEN_507;
  wire  GEN_259;
  reg [31:0] GEN_508;
  wire  GEN_260;
  reg [31:0] GEN_509;
  wire  GEN_261;
  reg [31:0] GEN_510;
  wire  GEN_262;
  reg [31:0] GEN_511;
  wire  GEN_263;
  reg [31:0] GEN_512;
  wire [2:0] GEN_264;
  reg [31:0] GEN_513;
  wire [1:0] GEN_265;
  reg [31:0] GEN_514;
  wire [64:0] GEN_266;
  reg [95:0] GEN_515;
  wire [64:0] GEN_267;
  reg [95:0] GEN_516;
  wire [64:0] GEN_268;
  reg [95:0] GEN_517;
  wire  GEN_269;
  reg [31:0] GEN_518;
  IBuf ibuf (
    .clk(ibuf_clk),
    .reset(ibuf_reset),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(ibuf_io_imem_valid),
    .io_imem_bits_btb_valid(ibuf_io_imem_bits_btb_valid),
    .io_imem_bits_btb_bits_taken(ibuf_io_imem_bits_btb_bits_taken),
    .io_imem_bits_btb_bits_mask(ibuf_io_imem_bits_btb_bits_mask),
    .io_imem_bits_btb_bits_bridx(ibuf_io_imem_bits_btb_bits_bridx),
    .io_imem_bits_btb_bits_target(ibuf_io_imem_bits_btb_bits_target),
    .io_imem_bits_btb_bits_entry(ibuf_io_imem_bits_btb_bits_entry),
    .io_imem_bits_btb_bits_bht_history(ibuf_io_imem_bits_btb_bits_bht_history),
    .io_imem_bits_btb_bits_bht_value(ibuf_io_imem_bits_btb_bits_bht_value),
    .io_imem_bits_pc(ibuf_io_imem_bits_pc),
    .io_imem_bits_data(ibuf_io_imem_bits_data),
    .io_imem_bits_mask(ibuf_io_imem_bits_mask),
    .io_imem_bits_xcpt_if(ibuf_io_imem_bits_xcpt_if),
    .io_imem_bits_replay(ibuf_io_imem_bits_replay),
    .io_kill(ibuf_io_kill),
    .io_pc(ibuf_io_pc),
    .io_btb_resp_taken(ibuf_io_btb_resp_taken),
    .io_btb_resp_mask(ibuf_io_btb_resp_mask),
    .io_btb_resp_bridx(ibuf_io_btb_resp_bridx),
    .io_btb_resp_target(ibuf_io_btb_resp_target),
    .io_btb_resp_entry(ibuf_io_btb_resp_entry),
    .io_btb_resp_bht_history(ibuf_io_btb_resp_bht_history),
    .io_btb_resp_bht_value(ibuf_io_btb_resp_bht_value),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_inst_0_bits_pf0(ibuf_io_inst_0_bits_pf0),
    .io_inst_0_bits_pf1(ibuf_io_inst_0_bits_pf1),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_btb_hit(ibuf_io_inst_0_bits_btb_hit),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_inst_rs3(ibuf_io_inst_0_bits_inst_rs3)
  );
  CSRFile csr (
    .clk(csr_clk),
    .reset(csr_reset),
    .io_prci_reset(csr_io_prci_reset),
    .io_prci_id(csr_io_prci_id),
    .io_prci_interrupts_meip(csr_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(csr_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(csr_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(csr_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(csr_io_prci_interrupts_msip),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_csr_stall(csr_io_csr_stall),
    .io_csr_xcpt(csr_io_csr_xcpt),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero3(csr_io_status_zero3),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_vm(csr_io_status_vm),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_pum(csr_io_status_pum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_asid(csr_io_ptbr_asid),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_badaddr(csr_io_badaddr),
    .io_fatc(csr_io_fatc),
    .io_time(csr_io_time),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_rocc_cmd_ready(csr_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(csr_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(csr_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(csr_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(csr_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(csr_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(csr_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(csr_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(csr_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(csr_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(csr_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(csr_io_rocc_cmd_bits_rs2),
    .io_rocc_cmd_bits_status_debug(csr_io_rocc_cmd_bits_status_debug),
    .io_rocc_cmd_bits_status_prv(csr_io_rocc_cmd_bits_status_prv),
    .io_rocc_cmd_bits_status_sd(csr_io_rocc_cmd_bits_status_sd),
    .io_rocc_cmd_bits_status_zero3(csr_io_rocc_cmd_bits_status_zero3),
    .io_rocc_cmd_bits_status_sd_rv32(csr_io_rocc_cmd_bits_status_sd_rv32),
    .io_rocc_cmd_bits_status_zero2(csr_io_rocc_cmd_bits_status_zero2),
    .io_rocc_cmd_bits_status_vm(csr_io_rocc_cmd_bits_status_vm),
    .io_rocc_cmd_bits_status_zero1(csr_io_rocc_cmd_bits_status_zero1),
    .io_rocc_cmd_bits_status_mxr(csr_io_rocc_cmd_bits_status_mxr),
    .io_rocc_cmd_bits_status_pum(csr_io_rocc_cmd_bits_status_pum),
    .io_rocc_cmd_bits_status_mprv(csr_io_rocc_cmd_bits_status_mprv),
    .io_rocc_cmd_bits_status_xs(csr_io_rocc_cmd_bits_status_xs),
    .io_rocc_cmd_bits_status_fs(csr_io_rocc_cmd_bits_status_fs),
    .io_rocc_cmd_bits_status_mpp(csr_io_rocc_cmd_bits_status_mpp),
    .io_rocc_cmd_bits_status_hpp(csr_io_rocc_cmd_bits_status_hpp),
    .io_rocc_cmd_bits_status_spp(csr_io_rocc_cmd_bits_status_spp),
    .io_rocc_cmd_bits_status_mpie(csr_io_rocc_cmd_bits_status_mpie),
    .io_rocc_cmd_bits_status_hpie(csr_io_rocc_cmd_bits_status_hpie),
    .io_rocc_cmd_bits_status_spie(csr_io_rocc_cmd_bits_status_spie),
    .io_rocc_cmd_bits_status_upie(csr_io_rocc_cmd_bits_status_upie),
    .io_rocc_cmd_bits_status_mie(csr_io_rocc_cmd_bits_status_mie),
    .io_rocc_cmd_bits_status_hie(csr_io_rocc_cmd_bits_status_hie),
    .io_rocc_cmd_bits_status_sie(csr_io_rocc_cmd_bits_status_sie),
    .io_rocc_cmd_bits_status_uie(csr_io_rocc_cmd_bits_status_uie),
    .io_rocc_resp_ready(csr_io_rocc_resp_ready),
    .io_rocc_resp_valid(csr_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(csr_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(csr_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(csr_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(csr_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(csr_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(csr_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(csr_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(csr_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(csr_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(csr_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(csr_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(csr_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(csr_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(csr_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(csr_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(csr_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(csr_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(csr_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(csr_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(csr_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(csr_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(csr_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(csr_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(csr_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(csr_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(csr_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(csr_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(csr_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(csr_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(csr_io_rocc_mem_ordered),
    .io_rocc_busy(csr_io_rocc_busy),
    .io_rocc_interrupt(csr_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(csr_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(csr_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(csr_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(csr_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(csr_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(csr_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(csr_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(csr_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(csr_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(csr_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(csr_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(csr_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(csr_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(csr_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(csr_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(csr_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(csr_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(csr_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(csr_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(csr_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(csr_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(csr_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(csr_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(csr_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(csr_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(csr_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(csr_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(csr_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(csr_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(csr_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(csr_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(csr_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(csr_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(csr_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(csr_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(csr_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(csr_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(csr_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(csr_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(csr_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(csr_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(csr_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(csr_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(csr_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(csr_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(csr_io_rocc_exception),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_ttype(csr_io_bp_0_control_ttype),
    .io_bp_0_control_dmode(csr_io_bp_0_control_dmode),
    .io_bp_0_control_maskmax(csr_io_bp_0_control_maskmax),
    .io_bp_0_control_reserved(csr_io_bp_0_control_reserved),
    .io_bp_0_control_action(csr_io_bp_0_control_action),
    .io_bp_0_control_chain(csr_io_bp_0_control_chain),
    .io_bp_0_control_zero(csr_io_bp_0_control_zero),
    .io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_h(csr_io_bp_0_control_h),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_address(csr_io_bp_0_address)
  );
  BreakpointUnit bpu (
    .clk(bpu_clk),
    .reset(bpu_reset),
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_status_sd(bpu_io_status_sd),
    .io_status_zero3(bpu_io_status_zero3),
    .io_status_sd_rv32(bpu_io_status_sd_rv32),
    .io_status_zero2(bpu_io_status_zero2),
    .io_status_vm(bpu_io_status_vm),
    .io_status_zero1(bpu_io_status_zero1),
    .io_status_mxr(bpu_io_status_mxr),
    .io_status_pum(bpu_io_status_pum),
    .io_status_mprv(bpu_io_status_mprv),
    .io_status_xs(bpu_io_status_xs),
    .io_status_fs(bpu_io_status_fs),
    .io_status_mpp(bpu_io_status_mpp),
    .io_status_hpp(bpu_io_status_hpp),
    .io_status_spp(bpu_io_status_spp),
    .io_status_mpie(bpu_io_status_mpie),
    .io_status_hpie(bpu_io_status_hpie),
    .io_status_spie(bpu_io_status_spie),
    .io_status_upie(bpu_io_status_upie),
    .io_status_mie(bpu_io_status_mie),
    .io_status_hie(bpu_io_status_hie),
    .io_status_sie(bpu_io_status_sie),
    .io_status_uie(bpu_io_status_uie),
    .io_bp_0_control_ttype(bpu_io_bp_0_control_ttype),
    .io_bp_0_control_dmode(bpu_io_bp_0_control_dmode),
    .io_bp_0_control_maskmax(bpu_io_bp_0_control_maskmax),
    .io_bp_0_control_reserved(bpu_io_bp_0_control_reserved),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_chain(bpu_io_bp_0_control_chain),
    .io_bp_0_control_zero(bpu_io_bp_0_control_zero),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_h(bpu_io_bp_0_control_h),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st),
    .io_debug_if(bpu_io_debug_if),
    .io_debug_ld(bpu_io_debug_ld),
    .io_debug_st(bpu_io_debug_st)
  );
  ALU alu (
    .clk(alu_clk),
    .reset(alu_reset),
    .io_dw(alu_io_dw),
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  MulDiv div (
    .clk(div_clk),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_dw(div_io_req_bits_dw),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag)
  );
  assign io_imem_req_valid = take_pc_mem_wb;
  assign io_imem_req_bits_pc = T_8120;
  assign io_imem_req_bits_speculative = T_7902;
  assign io_imem_resp_ready = ibuf_io_imem_ready;
  assign io_imem_btb_update_valid = T_8137;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign io_imem_btb_update_bits_pc = T_8156;
  assign io_imem_btb_update_bits_target = io_imem_req_bits_pc[38:0];
  assign io_imem_btb_update_bits_taken = GEN_155;
  assign io_imem_btb_update_bits_isValid = T_8140;
  assign io_imem_btb_update_bits_isJump = T_8141;
  assign io_imem_btb_update_bits_isReturn = T_8147;
  assign io_imem_btb_update_bits_br_pc = T_8152[38:0];
  assign io_imem_bht_update_valid = T_8160;
  assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_pc = io_imem_btb_update_bits_pc;
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_mispredict = mem_wrong_npc;
  assign io_imem_ras_update_valid = T_8131;
  assign io_imem_ras_update_bits_isCall = T_8165;
  assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
  assign io_imem_ras_update_bits_returnAddr = mem_int_wdata[38:0];
  assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_flush_icache = T_8124;
  assign io_imem_flush_tlb = csr_io_fatc;
  assign io_dmem_req_valid = T_8170;
  assign io_dmem_req_bits_addr = T_8195;
  assign io_dmem_req_bits_tag = ex_dcache_tag;
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_data = GEN_156;
  assign io_dmem_s1_kill = T_8197;
  assign io_dmem_s1_data = T_8196;
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_ptw_ptbr_asid = csr_io_ptbr_asid;
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn;
  assign io_ptw_invalidate = csr_io_fatc;
  assign io_ptw_status_debug = csr_io_status_debug;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_sd = csr_io_status_sd;
  assign io_ptw_status_zero3 = csr_io_status_zero3;
  assign io_ptw_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_ptw_status_zero2 = csr_io_status_zero2;
  assign io_ptw_status_vm = csr_io_status_vm;
  assign io_ptw_status_zero1 = csr_io_status_zero1;
  assign io_ptw_status_mxr = csr_io_status_mxr;
  assign io_ptw_status_pum = csr_io_status_pum;
  assign io_ptw_status_mprv = csr_io_status_mprv;
  assign io_ptw_status_xs = csr_io_status_xs;
  assign io_ptw_status_fs = csr_io_status_fs;
  assign io_ptw_status_mpp = csr_io_status_mpp;
  assign io_ptw_status_hpp = csr_io_status_hpp;
  assign io_ptw_status_spp = csr_io_status_spp;
  assign io_ptw_status_mpie = csr_io_status_mpie;
  assign io_ptw_status_hpie = csr_io_status_hpie;
  assign io_ptw_status_spie = csr_io_status_spie;
  assign io_ptw_status_upie = csr_io_status_upie;
  assign io_ptw_status_mie = csr_io_status_mie;
  assign io_ptw_status_hie = csr_io_status_hie;
  assign io_ptw_status_sie = csr_io_status_sie;
  assign io_ptw_status_uie = csr_io_status_uie;
  assign io_fpu_inst = ibuf_io_inst_0_bits_inst_bits;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_dmem_resp_val = T_8169;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_tag = dmem_resp_waddr;
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass;
  assign io_fpu_valid = T_8168;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_killm = killm_common;
  assign io_fpu_cp_req_valid = GEN_157;
  assign io_fpu_cp_req_bits_cmd = GEN_158;
  assign io_fpu_cp_req_bits_ldst = GEN_159;
  assign io_fpu_cp_req_bits_wen = GEN_162;
  assign io_fpu_cp_req_bits_ren1 = GEN_163;
  assign io_fpu_cp_req_bits_ren2 = GEN_165;
  assign io_fpu_cp_req_bits_ren3 = GEN_166;
  assign io_fpu_cp_req_bits_swap12 = GEN_174;
  assign io_fpu_cp_req_bits_swap23 = GEN_175;
  assign io_fpu_cp_req_bits_single = GEN_176;
  assign io_fpu_cp_req_bits_fromint = GEN_177;
  assign io_fpu_cp_req_bits_toint = GEN_178;
  assign io_fpu_cp_req_bits_fastpipe = GEN_179;
  assign io_fpu_cp_req_bits_fma = GEN_180;
  assign io_fpu_cp_req_bits_div = GEN_181;
  assign io_fpu_cp_req_bits_sqrt = GEN_182;
  assign io_fpu_cp_req_bits_round = GEN_183;
  assign io_fpu_cp_req_bits_wflags = GEN_184;
  assign io_fpu_cp_req_bits_rm = GEN_185;
  assign io_fpu_cp_req_bits_typ = GEN_186;
  assign io_fpu_cp_req_bits_in1 = GEN_187;
  assign io_fpu_cp_req_bits_in2 = GEN_188;
  assign io_fpu_cp_req_bits_in3 = GEN_189;
  assign io_fpu_cp_resp_ready = GEN_190;
  assign io_rocc_cmd_valid = T_8212;
  assign io_rocc_cmd_bits_inst_funct = T_8234_funct;
  assign io_rocc_cmd_bits_inst_rs2 = T_8234_rs2;
  assign io_rocc_cmd_bits_inst_rs1 = T_8234_rs1;
  assign io_rocc_cmd_bits_inst_xd = T_8234_xd;
  assign io_rocc_cmd_bits_inst_xs1 = T_8234_xs1;
  assign io_rocc_cmd_bits_inst_xs2 = T_8234_xs2;
  assign io_rocc_cmd_bits_inst_rd = T_8234_rd;
  assign io_rocc_cmd_bits_inst_opcode = T_8234_opcode;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign io_rocc_cmd_bits_status_debug = csr_io_status_debug;
  assign io_rocc_cmd_bits_status_prv = csr_io_status_prv;
  assign io_rocc_cmd_bits_status_sd = csr_io_status_sd;
  assign io_rocc_cmd_bits_status_zero3 = csr_io_status_zero3;
  assign io_rocc_cmd_bits_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_rocc_cmd_bits_status_zero2 = csr_io_status_zero2;
  assign io_rocc_cmd_bits_status_vm = csr_io_status_vm;
  assign io_rocc_cmd_bits_status_zero1 = csr_io_status_zero1;
  assign io_rocc_cmd_bits_status_mxr = csr_io_status_mxr;
  assign io_rocc_cmd_bits_status_pum = csr_io_status_pum;
  assign io_rocc_cmd_bits_status_mprv = csr_io_status_mprv;
  assign io_rocc_cmd_bits_status_xs = csr_io_status_xs;
  assign io_rocc_cmd_bits_status_fs = csr_io_status_fs;
  assign io_rocc_cmd_bits_status_mpp = csr_io_status_mpp;
  assign io_rocc_cmd_bits_status_hpp = csr_io_status_hpp;
  assign io_rocc_cmd_bits_status_spp = csr_io_status_spp;
  assign io_rocc_cmd_bits_status_mpie = csr_io_status_mpie;
  assign io_rocc_cmd_bits_status_hpie = csr_io_status_hpie;
  assign io_rocc_cmd_bits_status_spie = csr_io_status_spie;
  assign io_rocc_cmd_bits_status_upie = csr_io_status_upie;
  assign io_rocc_cmd_bits_status_mie = csr_io_status_mie;
  assign io_rocc_cmd_bits_status_hie = csr_io_status_hie;
  assign io_rocc_cmd_bits_status_sie = csr_io_status_sie;
  assign io_rocc_cmd_bits_status_uie = csr_io_status_uie;
  assign io_rocc_resp_ready = GEN_191;
  assign io_rocc_mem_req_ready = GEN_192;
  assign io_rocc_mem_s2_nack = GEN_193;
  assign io_rocc_mem_resp_valid = GEN_194;
  assign io_rocc_mem_resp_bits_addr = GEN_195;
  assign io_rocc_mem_resp_bits_tag = GEN_196;
  assign io_rocc_mem_resp_bits_cmd = GEN_197;
  assign io_rocc_mem_resp_bits_typ = GEN_198;
  assign io_rocc_mem_resp_bits_data = GEN_199;
  assign io_rocc_mem_resp_bits_replay = GEN_200;
  assign io_rocc_mem_resp_bits_has_data = GEN_201;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_202;
  assign io_rocc_mem_resp_bits_store_data = GEN_203;
  assign io_rocc_mem_replay_next = GEN_204;
  assign io_rocc_mem_xcpt_ma_ld = GEN_205;
  assign io_rocc_mem_xcpt_ma_st = GEN_206;
  assign io_rocc_mem_xcpt_pf_ld = GEN_207;
  assign io_rocc_mem_xcpt_pf_st = GEN_208;
  assign io_rocc_mem_ordered = GEN_209;
  assign io_rocc_autl_acquire_ready = GEN_210;
  assign io_rocc_autl_grant_valid = GEN_211;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_212;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_213;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_214;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_215;
  assign io_rocc_autl_grant_bits_g_type = GEN_216;
  assign io_rocc_autl_grant_bits_data = GEN_217;
  assign io_rocc_fpu_req_ready = GEN_218;
  assign io_rocc_fpu_resp_valid = GEN_219;
  assign io_rocc_fpu_resp_bits_data = GEN_220;
  assign io_rocc_fpu_resp_bits_exc = GEN_221;
  assign io_rocc_exception = T_8215;
  assign take_pc_mem = T_7829;
  assign take_pc_wb = T_7919;
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem;
  assign ibuf_clk = clk;
  assign ibuf_reset = reset;
  assign ibuf_io_imem_valid = io_imem_resp_valid;
  assign ibuf_io_imem_bits_btb_valid = io_imem_resp_bits_btb_valid;
  assign ibuf_io_imem_bits_btb_bits_taken = io_imem_resp_bits_btb_bits_taken;
  assign ibuf_io_imem_bits_btb_bits_mask = io_imem_resp_bits_btb_bits_mask;
  assign ibuf_io_imem_bits_btb_bits_bridx = io_imem_resp_bits_btb_bits_bridx;
  assign ibuf_io_imem_bits_btb_bits_target = io_imem_resp_bits_btb_bits_target;
  assign ibuf_io_imem_bits_btb_bits_entry = io_imem_resp_bits_btb_bits_entry;
  assign ibuf_io_imem_bits_btb_bits_bht_history = io_imem_resp_bits_btb_bits_bht_history;
  assign ibuf_io_imem_bits_btb_bits_bht_value = io_imem_resp_bits_btb_bits_bht_value;
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc;
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data;
  assign ibuf_io_imem_bits_mask = io_imem_resp_bits_mask;
  assign ibuf_io_imem_bits_xcpt_if = io_imem_resp_bits_xcpt_if;
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay;
  assign ibuf_io_kill = take_pc_mem_wb;
  assign ibuf_io_inst_0_ready = T_8127;
  assign id_ctrl_legal = T_6778;
  assign id_ctrl_fp = 1'h0;
  assign id_ctrl_rocc = 1'h0;
  assign id_ctrl_branch = T_6784;
  assign id_ctrl_jal = T_6790;
  assign id_ctrl_jalr = T_6796;
  assign id_ctrl_rxs2 = T_6814;
  assign id_ctrl_rxs1 = T_6835;
  assign id_ctrl_sel_alu2 = T_6871;
  assign id_ctrl_sel_alu1 = T_6888;
  assign id_ctrl_sel_imm = T_6920;
  assign id_ctrl_alu_dw = T_6931;
  assign id_ctrl_alu_fn = T_7015;
  assign id_ctrl_mem = T_7031;
  assign id_ctrl_mem_cmd = T_7091;
  assign id_ctrl_mem_type = T_7111;
  assign id_ctrl_rfs1 = 1'h0;
  assign id_ctrl_rfs2 = 1'h0;
  assign id_ctrl_rfs3 = 1'h0;
  assign id_ctrl_wfd = 1'h0;
  assign id_ctrl_div = T_7119;
  assign id_ctrl_wxd = T_7149;
  assign id_ctrl_csr = T_7169;
  assign id_ctrl_fence_i = T_7173;
  assign id_ctrl_fence = T_7179;
  assign id_ctrl_amo = T_7185;
  assign T_6645 = ibuf_io_inst_0_bits_inst_bits & 32'h405f;
  assign T_6647 = T_6645 == 32'h3;
  assign T_6649 = ibuf_io_inst_0_bits_inst_bits & 32'h207f;
  assign T_6651 = T_6649 == 32'h3;
  assign T_6653 = ibuf_io_inst_0_bits_inst_bits & 32'h106f;
  assign T_6655 = T_6653 == 32'h3;
  assign T_6657 = ibuf_io_inst_0_bits_inst_bits & 32'h607f;
  assign T_6659 = T_6657 == 32'hf;
  assign T_6661 = ibuf_io_inst_0_bits_inst_bits & 32'h7077;
  assign T_6663 = T_6661 == 32'h13;
  assign T_6665 = ibuf_io_inst_0_bits_inst_bits & 32'h5f;
  assign T_6667 = T_6665 == 32'h17;
  assign T_6669 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00007f;
  assign T_6671 = T_6669 == 32'h33;
  assign T_6673 = ibuf_io_inst_0_bits_inst_bits & 32'hbe007077;
  assign T_6675 = T_6673 == 32'h33;
  assign T_6677 = ibuf_io_inst_0_bits_inst_bits & 32'h707b;
  assign T_6679 = T_6677 == 32'h63;
  assign T_6681 = ibuf_io_inst_0_bits_inst_bits & 32'h7f;
  assign T_6683 = T_6681 == 32'h6f;
  assign T_6685 = ibuf_io_inst_0_bits_inst_bits & 32'hffefffff;
  assign T_6687 = T_6685 == 32'h73;
  assign T_6689 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00305f;
  assign T_6691 = T_6689 == 32'h1013;
  assign T_6693 = ibuf_io_inst_0_bits_inst_bits & 32'hfe00305f;
  assign T_6695 = T_6693 == 32'h101b;
  assign T_6699 = T_6649 == 32'h2013;
  assign T_6701 = ibuf_io_inst_0_bits_inst_bits & 32'h1800607f;
  assign T_6703 = T_6701 == 32'h202f;
  assign T_6707 = T_6649 == 32'h2073;
  assign T_6709 = ibuf_io_inst_0_bits_inst_bits & 32'hbc00707f;
  assign T_6711 = T_6709 == 32'h5013;
  assign T_6713 = ibuf_io_inst_0_bits_inst_bits & 32'hbe00705f;
  assign T_6715 = T_6713 == 32'h501b;
  assign T_6719 = T_6673 == 32'h5033;
  assign T_6721 = ibuf_io_inst_0_bits_inst_bits & 32'hfe004077;
  assign T_6723 = T_6721 == 32'h2004033;
  assign T_6725 = ibuf_io_inst_0_bits_inst_bits & 32'he800607f;
  assign T_6727 = T_6725 == 32'h800202f;
  assign T_6729 = ibuf_io_inst_0_bits_inst_bits & 32'hf9f0607f;
  assign T_6731 = T_6729 == 32'h1000202f;
  assign T_6733 = ibuf_io_inst_0_bits_inst_bits == 32'h10500073;
  assign T_6735 = ibuf_io_inst_0_bits_inst_bits == 32'h30200073;
  assign T_6737 = ibuf_io_inst_0_bits_inst_bits == 32'h7b200073;
  assign T_6739 = ibuf_io_inst_0_bits_inst_bits & 32'h306f;
  assign T_6741 = T_6739 == 32'h1063;
  assign T_6743 = ibuf_io_inst_0_bits_inst_bits & 32'h407f;
  assign T_6745 = T_6743 == 32'h4063;
  assign T_6747 = ibuf_io_inst_0_bits_inst_bits & 32'hfc007077;
  assign T_6749 = T_6747 == 32'h33;
  assign T_6752 = T_6647 | T_6651;
  assign T_6753 = T_6752 | T_6655;
  assign T_6754 = T_6753 | T_6659;
  assign T_6755 = T_6754 | T_6663;
  assign T_6756 = T_6755 | T_6667;
  assign T_6757 = T_6756 | T_6671;
  assign T_6758 = T_6757 | T_6675;
  assign T_6759 = T_6758 | T_6679;
  assign T_6760 = T_6759 | T_6683;
  assign T_6761 = T_6760 | T_6687;
  assign T_6762 = T_6761 | T_6691;
  assign T_6763 = T_6762 | T_6695;
  assign T_6764 = T_6763 | T_6699;
  assign T_6765 = T_6764 | T_6703;
  assign T_6766 = T_6765 | T_6707;
  assign T_6767 = T_6766 | T_6711;
  assign T_6768 = T_6767 | T_6715;
  assign T_6769 = T_6768 | T_6719;
  assign T_6770 = T_6769 | T_6723;
  assign T_6771 = T_6770 | T_6727;
  assign T_6772 = T_6771 | T_6731;
  assign T_6773 = T_6772 | T_6733;
  assign T_6774 = T_6773 | T_6735;
  assign T_6775 = T_6774 | T_6737;
  assign T_6776 = T_6775 | T_6741;
  assign T_6777 = T_6776 | T_6745;
  assign T_6778 = T_6777 | T_6749;
  assign T_6782 = ibuf_io_inst_0_bits_inst_bits & 32'h54;
  assign T_6784 = T_6782 == 32'h40;
  assign T_6788 = ibuf_io_inst_0_bits_inst_bits & 32'h48;
  assign T_6790 = T_6788 == 32'h48;
  assign T_6794 = ibuf_io_inst_0_bits_inst_bits & 32'h1c;
  assign T_6796 = T_6794 == 32'h4;
  assign T_6800 = ibuf_io_inst_0_bits_inst_bits & 32'h70;
  assign T_6802 = T_6800 == 32'h20;
  assign T_6804 = ibuf_io_inst_0_bits_inst_bits & 32'h64;
  assign T_6806 = T_6804 == 32'h20;
  assign T_6808 = ibuf_io_inst_0_bits_inst_bits & 32'h34;
  assign T_6810 = T_6808 == 32'h20;
  assign T_6813 = T_6802 | T_6806;
  assign T_6814 = T_6813 | T_6810;
  assign T_6816 = ibuf_io_inst_0_bits_inst_bits & 32'h4004;
  assign T_6818 = T_6816 == 32'h0;
  assign T_6820 = ibuf_io_inst_0_bits_inst_bits & 32'h44;
  assign T_6822 = T_6820 == 32'h0;
  assign T_6824 = ibuf_io_inst_0_bits_inst_bits & 32'h18;
  assign T_6826 = T_6824 == 32'h0;
  assign T_6828 = ibuf_io_inst_0_bits_inst_bits & 32'h2050;
  assign T_6830 = T_6828 == 32'h2000;
  assign T_6833 = T_6818 | T_6822;
  assign T_6834 = T_6833 | T_6826;
  assign T_6835 = T_6834 | T_6830;
  assign T_6837 = ibuf_io_inst_0_bits_inst_bits & 32'h58;
  assign T_6839 = T_6837 == 32'h0;
  assign T_6841 = ibuf_io_inst_0_bits_inst_bits & 32'h20;
  assign T_6843 = T_6841 == 32'h0;
  assign T_6845 = ibuf_io_inst_0_bits_inst_bits & 32'hc;
  assign T_6847 = T_6845 == 32'h4;
  assign T_6849 = ibuf_io_inst_0_bits_inst_bits & 32'h4050;
  assign T_6851 = T_6849 == 32'h4050;
  assign T_6854 = T_6839 | T_6843;
  assign T_6855 = T_6854 | T_6847;
  assign T_6856 = T_6855 | T_6790;
  assign T_6857 = T_6856 | T_6851;
  assign T_6861 = T_6788 == 32'h0;
  assign T_6863 = ibuf_io_inst_0_bits_inst_bits & 32'h4008;
  assign T_6865 = T_6863 == 32'h4000;
  assign T_6868 = T_6861 | T_6822;
  assign T_6869 = T_6868 | T_6826;
  assign T_6870 = T_6869 | T_6865;
  assign T_6871 = {T_6870,T_6857};
  assign T_6873 = ibuf_io_inst_0_bits_inst_bits & 32'h50;
  assign T_6875 = T_6873 == 32'h0;
  assign T_6878 = T_6818 | T_6875;
  assign T_6879 = T_6878 | T_6822;
  assign T_6880 = T_6879 | T_6826;
  assign T_6882 = ibuf_io_inst_0_bits_inst_bits & 32'h24;
  assign T_6884 = T_6882 == 32'h4;
  assign T_6887 = T_6884 | T_6790;
  assign T_6888 = {T_6887,T_6880};
  assign T_6892 = T_6824 == 32'h8;
  assign T_6896 = T_6820 == 32'h40;
  assign T_6899 = T_6892 | T_6896;
  assign T_6903 = T_6820 == 32'h4;
  assign T_6906 = T_6903 | T_6892;
  assign T_6910 = T_6882 == 32'h0;
  assign T_6912 = ibuf_io_inst_0_bits_inst_bits & 32'h14;
  assign T_6914 = T_6912 == 32'h10;
  assign T_6917 = T_6910 | T_6796;
  assign T_6918 = T_6917 | T_6914;
  assign T_6919 = {T_6918,T_6906};
  assign T_6920 = {T_6919,T_6899};
  assign T_6922 = ibuf_io_inst_0_bits_inst_bits & 32'h10;
  assign T_6924 = T_6922 == 32'h0;
  assign T_6926 = ibuf_io_inst_0_bits_inst_bits & 32'h8;
  assign T_6928 = T_6926 == 32'h0;
  assign T_6931 = T_6924 | T_6928;
  assign T_6933 = ibuf_io_inst_0_bits_inst_bits & 32'h3054;
  assign T_6935 = T_6933 == 32'h1010;
  assign T_6937 = ibuf_io_inst_0_bits_inst_bits & 32'h1058;
  assign T_6939 = T_6937 == 32'h1040;
  assign T_6941 = ibuf_io_inst_0_bits_inst_bits & 32'h7044;
  assign T_6943 = T_6941 == 32'h7000;
  assign T_6946 = T_6935 | T_6939;
  assign T_6947 = T_6946 | T_6943;
  assign T_6949 = ibuf_io_inst_0_bits_inst_bits & 32'h4054;
  assign T_6951 = T_6949 == 32'h40;
  assign T_6953 = ibuf_io_inst_0_bits_inst_bits & 32'h2058;
  assign T_6955 = T_6953 == 32'h2040;
  assign T_6959 = T_6933 == 32'h3010;
  assign T_6961 = ibuf_io_inst_0_bits_inst_bits & 32'h6054;
  assign T_6963 = T_6961 == 32'h6010;
  assign T_6965 = ibuf_io_inst_0_bits_inst_bits & 32'h40003034;
  assign T_6967 = T_6965 == 32'h40000030;
  assign T_6969 = ibuf_io_inst_0_bits_inst_bits & 32'h40001054;
  assign T_6971 = T_6969 == 32'h40001010;
  assign T_6974 = T_6951 | T_6955;
  assign T_6975 = T_6974 | T_6959;
  assign T_6976 = T_6975 | T_6963;
  assign T_6977 = T_6976 | T_6967;
  assign T_6978 = T_6977 | T_6971;
  assign T_6980 = ibuf_io_inst_0_bits_inst_bits & 32'h2054;
  assign T_6982 = T_6980 == 32'h2010;
  assign T_6984 = ibuf_io_inst_0_bits_inst_bits & 32'h40004054;
  assign T_6986 = T_6984 == 32'h4010;
  assign T_6988 = ibuf_io_inst_0_bits_inst_bits & 32'h5054;
  assign T_6990 = T_6988 == 32'h4010;
  assign T_6992 = ibuf_io_inst_0_bits_inst_bits & 32'h4058;
  assign T_6994 = T_6992 == 32'h4040;
  assign T_6997 = T_6982 | T_6986;
  assign T_6998 = T_6997 | T_6990;
  assign T_6999 = T_6998 | T_6994;
  assign T_7003 = T_6961 == 32'h2010;
  assign T_7005 = ibuf_io_inst_0_bits_inst_bits & 32'h40003054;
  assign T_7007 = T_7005 == 32'h40001010;
  assign T_7010 = T_7003 | T_6994;
  assign T_7011 = T_7010 | T_6967;
  assign T_7012 = T_7011 | T_7007;
  assign T_7013 = {T_6978,T_6947};
  assign T_7014 = {T_7012,T_6999};
  assign T_7015 = {T_7014,T_7013};
  assign T_7017 = ibuf_io_inst_0_bits_inst_bits & 32'h107f;
  assign T_7019 = T_7017 == 32'h3;
  assign T_7021 = ibuf_io_inst_0_bits_inst_bits & 32'h707f;
  assign T_7023 = T_7021 == 32'h100f;
  assign T_7027 = T_6752 | T_7019;
  assign T_7028 = T_7027 | T_7023;
  assign T_7029 = T_7028 | T_6703;
  assign T_7030 = T_7029 | T_6727;
  assign T_7031 = T_7030 | T_6731;
  assign T_7033 = ibuf_io_inst_0_bits_inst_bits & 32'h2008;
  assign T_7035 = T_7033 == 32'h8;
  assign T_7037 = ibuf_io_inst_0_bits_inst_bits & 32'h28;
  assign T_7039 = T_7037 == 32'h20;
  assign T_7041 = ibuf_io_inst_0_bits_inst_bits & 32'h18000020;
  assign T_7043 = T_7041 == 32'h18000020;
  assign T_7045 = ibuf_io_inst_0_bits_inst_bits & 32'h20000020;
  assign T_7047 = T_7045 == 32'h20000020;
  assign T_7050 = T_7035 | T_7039;
  assign T_7051 = T_7050 | T_7043;
  assign T_7052 = T_7051 | T_7047;
  assign T_7054 = ibuf_io_inst_0_bits_inst_bits & 32'h10002008;
  assign T_7056 = T_7054 == 32'h10002008;
  assign T_7058 = ibuf_io_inst_0_bits_inst_bits & 32'h40002008;
  assign T_7060 = T_7058 == 32'h40002008;
  assign T_7063 = T_7056 | T_7060;
  assign T_7065 = ibuf_io_inst_0_bits_inst_bits & 32'h8000008;
  assign T_7067 = T_7065 == 32'h8000008;
  assign T_7069 = ibuf_io_inst_0_bits_inst_bits & 32'h10000008;
  assign T_7071 = T_7069 == 32'h10000008;
  assign T_7073 = ibuf_io_inst_0_bits_inst_bits & 32'h80000008;
  assign T_7075 = T_7073 == 32'h80000008;
  assign T_7078 = T_7035 | T_7067;
  assign T_7079 = T_7078 | T_7071;
  assign T_7080 = T_7079 | T_7075;
  assign T_7082 = ibuf_io_inst_0_bits_inst_bits & 32'h18002008;
  assign T_7084 = T_7082 == 32'h2008;
  assign T_7088 = {T_7063,T_7052};
  assign T_7089 = {1'h0,T_7084};
  assign T_7090 = {T_7089,T_7080};
  assign T_7091 = {T_7090,T_7088};
  assign T_7093 = ibuf_io_inst_0_bits_inst_bits & 32'h1000;
  assign T_7095 = T_7093 == 32'h1000;
  assign T_7099 = ibuf_io_inst_0_bits_inst_bits & 32'h2000;
  assign T_7101 = T_7099 == 32'h2000;
  assign T_7105 = ibuf_io_inst_0_bits_inst_bits & 32'h4000;
  assign T_7107 = T_7105 == 32'h4000;
  assign T_7110 = {T_7107,T_7101};
  assign T_7111 = {T_7110,T_7095};
  assign T_7117 = ibuf_io_inst_0_bits_inst_bits & 32'h2000074;
  assign T_7119 = T_7117 == 32'h2000030;
  assign T_7125 = T_6873 == 32'h10;
  assign T_7127 = ibuf_io_inst_0_bits_inst_bits & 32'h1010;
  assign T_7129 = T_7127 == 32'h1010;
  assign T_7133 = T_7033 == 32'h2008;
  assign T_7135 = ibuf_io_inst_0_bits_inst_bits & 32'h2010;
  assign T_7137 = T_7135 == 32'h2010;
  assign T_7141 = T_7037 == 32'h0;
  assign T_7144 = T_6847 | T_7125;
  assign T_7145 = T_7144 | T_6790;
  assign T_7146 = T_7145 | T_7129;
  assign T_7147 = T_7146 | T_7133;
  assign T_7148 = T_7147 | T_7137;
  assign T_7149 = T_7148 | T_7141;
  assign T_7151 = ibuf_io_inst_0_bits_inst_bits & 32'h1050;
  assign T_7153 = T_7151 == 32'h1050;
  assign T_7159 = T_6828 == 32'h2050;
  assign T_7163 = ibuf_io_inst_0_bits_inst_bits & 32'h3050;
  assign T_7165 = T_7163 == 32'h50;
  assign T_7168 = {T_7165,T_7159};
  assign T_7169 = {T_7168,T_7153};
  assign T_7171 = ibuf_io_inst_0_bits_inst_bits & 32'h3058;
  assign T_7173 = T_7171 == 32'h1008;
  assign T_7179 = T_7171 == 32'h8;
  assign T_7183 = ibuf_io_inst_0_bits_inst_bits & 32'h6048;
  assign T_7185 = T_7183 == 32'h2008;
  assign id_load_use = T_8065;
  assign T_7192_T_7201_addr = T_7200;
  assign T_7192_T_7201_en = 1'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_7192_T_7201_data = T_7192[T_7192_T_7201_addr];
  `else
  assign T_7192_T_7201_data = T_7192_T_7201_addr >= 5'h1f ? GEN_398[63:0] : T_7192[T_7192_T_7201_addr];
  `endif
  assign T_7192_T_7211_addr = T_7210;
  assign T_7192_T_7211_en = 1'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_7192_T_7211_data = T_7192[T_7192_T_7211_addr];
  `else
  assign T_7192_T_7211_data = T_7192_T_7211_addr >= 5'h1f ? GEN_399[63:0] : T_7192[T_7192_T_7211_addr];
  `endif
  assign T_7192_T_7944_data = rf_wdata;
  assign T_7192_T_7944_addr = T_7943;
  assign T_7192_T_7944_mask = GEN_164;
  assign T_7192_T_7944_en = GEN_164;
  assign id_rs_0 = GEN_167;
  assign T_7196 = ibuf_io_inst_0_bits_inst_rs1 == 5'h0;
  assign T_7199 = ibuf_io_inst_0_bits_inst_rs1;
  assign T_7200 = ~ T_7199;
  assign T_7202 = T_7192_T_7201_data;
  assign id_rs_1 = GEN_168;
  assign T_7209 = ibuf_io_inst_0_bits_inst_rs2;
  assign T_7210 = ~ T_7209;
  assign T_7212 = T_7192_T_7211_data;
  assign ctrl_killd = T_8115;
  assign csr_clk = clk;
  assign csr_reset = reset;
  assign csr_io_prci_reset = io_prci_reset;
  assign csr_io_prci_id = io_prci_id;
  assign csr_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign csr_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign csr_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign csr_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign csr_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign csr_io_rw_addr = T_7971;
  assign csr_io_rw_cmd = T_7972;
  assign csr_io_rw_wdata = wb_reg_wdata;
  assign csr_io_exception = wb_reg_xcpt;
  assign csr_io_retire = wb_valid;
  assign csr_io_cause = wb_reg_cause;
  assign csr_io_pc = wb_reg_pc;
  assign csr_io_badaddr = T_7970;
  assign csr_io_fcsr_flags_valid = io_fpu_fcsr_flags_valid;
  assign csr_io_fcsr_flags_bits = io_fpu_fcsr_flags_bits;
  assign csr_io_rocc_cmd_ready = GEN_222;
  assign csr_io_rocc_resp_valid = GEN_223;
  assign csr_io_rocc_resp_bits_rd = GEN_224;
  assign csr_io_rocc_resp_bits_data = GEN_225;
  assign csr_io_rocc_mem_req_valid = GEN_226;
  assign csr_io_rocc_mem_req_bits_addr = GEN_227;
  assign csr_io_rocc_mem_req_bits_tag = GEN_228;
  assign csr_io_rocc_mem_req_bits_cmd = GEN_229;
  assign csr_io_rocc_mem_req_bits_typ = GEN_230;
  assign csr_io_rocc_mem_req_bits_phys = GEN_231;
  assign csr_io_rocc_mem_req_bits_data = GEN_232;
  assign csr_io_rocc_mem_s1_kill = GEN_233;
  assign csr_io_rocc_mem_s1_data = GEN_234;
  assign csr_io_rocc_mem_invalidate_lr = GEN_235;
  assign csr_io_rocc_busy = GEN_236;
  assign csr_io_rocc_interrupt = io_rocc_interrupt;
  assign csr_io_rocc_autl_acquire_valid = GEN_237;
  assign csr_io_rocc_autl_acquire_bits_addr_block = GEN_238;
  assign csr_io_rocc_autl_acquire_bits_client_xact_id = GEN_239;
  assign csr_io_rocc_autl_acquire_bits_addr_beat = GEN_240;
  assign csr_io_rocc_autl_acquire_bits_is_builtin_type = GEN_241;
  assign csr_io_rocc_autl_acquire_bits_a_type = GEN_242;
  assign csr_io_rocc_autl_acquire_bits_union = GEN_243;
  assign csr_io_rocc_autl_acquire_bits_data = GEN_244;
  assign csr_io_rocc_autl_grant_ready = GEN_245;
  assign csr_io_rocc_fpu_req_valid = GEN_246;
  assign csr_io_rocc_fpu_req_bits_cmd = GEN_247;
  assign csr_io_rocc_fpu_req_bits_ldst = GEN_248;
  assign csr_io_rocc_fpu_req_bits_wen = GEN_249;
  assign csr_io_rocc_fpu_req_bits_ren1 = GEN_250;
  assign csr_io_rocc_fpu_req_bits_ren2 = GEN_251;
  assign csr_io_rocc_fpu_req_bits_ren3 = GEN_252;
  assign csr_io_rocc_fpu_req_bits_swap12 = GEN_253;
  assign csr_io_rocc_fpu_req_bits_swap23 = GEN_254;
  assign csr_io_rocc_fpu_req_bits_single = GEN_255;
  assign csr_io_rocc_fpu_req_bits_fromint = GEN_256;
  assign csr_io_rocc_fpu_req_bits_toint = GEN_257;
  assign csr_io_rocc_fpu_req_bits_fastpipe = GEN_258;
  assign csr_io_rocc_fpu_req_bits_fma = GEN_259;
  assign csr_io_rocc_fpu_req_bits_div = GEN_260;
  assign csr_io_rocc_fpu_req_bits_sqrt = GEN_261;
  assign csr_io_rocc_fpu_req_bits_round = GEN_262;
  assign csr_io_rocc_fpu_req_bits_wflags = GEN_263;
  assign csr_io_rocc_fpu_req_bits_rm = GEN_264;
  assign csr_io_rocc_fpu_req_bits_typ = GEN_265;
  assign csr_io_rocc_fpu_req_bits_in1 = GEN_266;
  assign csr_io_rocc_fpu_req_bits_in2 = GEN_267;
  assign csr_io_rocc_fpu_req_bits_in3 = GEN_268;
  assign csr_io_rocc_fpu_resp_ready = GEN_269;
  assign id_csr_en = id_ctrl_csr != 3'h0;
  assign id_system_insn = id_ctrl_csr == 3'h4;
  assign T_7214 = id_ctrl_csr == 3'h2;
  assign T_7215 = id_ctrl_csr == 3'h3;
  assign T_7216 = T_7214 | T_7215;
  assign id_csr_ren = T_7216 & T_7196;
  assign id_csr = id_csr_ren ? 3'h5 : id_ctrl_csr;
  assign id_csr_addr = ibuf_io_inst_0_bits_inst_bits[31:20];
  assign T_7220 = id_csr_ren == 1'h0;
  assign T_7221 = id_csr_en & T_7220;
  assign T_7351 = id_csr_addr & 12'h46;
  assign T_7353 = T_7351 == 12'h40;
  assign T_7355 = id_csr_addr & 12'h244;
  assign T_7357 = T_7355 == 12'h240;
  assign T_7360 = T_7353 | T_7357;
  assign T_7363 = T_7360 == 1'h0;
  assign T_7364 = T_7221 & T_7363;
  assign id_csr_flush = id_system_insn | T_7364;
  assign T_7366 = id_ctrl_legal == 1'h0;
  assign T_7368 = csr_io_status_fs != 2'h0;
  assign T_7370 = T_7368 == 1'h0;
  assign T_7371 = id_ctrl_fp & T_7370;
  assign T_7372 = T_7366 | T_7371;
  assign T_7374 = csr_io_status_xs != 2'h0;
  assign T_7376 = T_7374 == 1'h0;
  assign T_7377 = id_ctrl_rocc & T_7376;
  assign id_illegal_insn = T_7372 | T_7377;
  assign id_amo_aq = ibuf_io_inst_0_bits_inst_bits[26];
  assign id_amo_rl = ibuf_io_inst_0_bits_inst_bits[25];
  assign T_7378 = id_ctrl_amo & id_amo_rl;
  assign id_fence_next = id_ctrl_fence | T_7378;
  assign T_7380 = io_dmem_ordered == 1'h0;
  assign id_mem_busy = T_7380 | io_dmem_req_valid;
  assign T_7386 = wb_reg_valid & wb_ctrl_rocc;
  assign T_7388 = id_reg_fence & id_mem_busy;
  assign T_7389 = id_fence_next | T_7388;
  assign T_7391 = id_ctrl_amo & id_amo_aq;
  assign T_7392 = T_7391 | id_ctrl_fence_i;
  assign T_7393 = id_ctrl_mem | id_ctrl_rocc;
  assign T_7394 = id_reg_fence & T_7393;
  assign T_7395 = T_7392 | T_7394;
  assign T_7396 = T_7395 | id_csr_en;
  assign T_7397 = id_mem_busy & T_7396;
  assign bpu_clk = clk;
  assign bpu_reset = reset;
  assign bpu_io_status_debug = csr_io_status_debug;
  assign bpu_io_status_prv = csr_io_status_prv;
  assign bpu_io_status_sd = csr_io_status_sd;
  assign bpu_io_status_zero3 = csr_io_status_zero3;
  assign bpu_io_status_sd_rv32 = csr_io_status_sd_rv32;
  assign bpu_io_status_zero2 = csr_io_status_zero2;
  assign bpu_io_status_vm = csr_io_status_vm;
  assign bpu_io_status_zero1 = csr_io_status_zero1;
  assign bpu_io_status_mxr = csr_io_status_mxr;
  assign bpu_io_status_pum = csr_io_status_pum;
  assign bpu_io_status_mprv = csr_io_status_mprv;
  assign bpu_io_status_xs = csr_io_status_xs;
  assign bpu_io_status_fs = csr_io_status_fs;
  assign bpu_io_status_mpp = csr_io_status_mpp;
  assign bpu_io_status_hpp = csr_io_status_hpp;
  assign bpu_io_status_spp = csr_io_status_spp;
  assign bpu_io_status_mpie = csr_io_status_mpie;
  assign bpu_io_status_hpie = csr_io_status_hpie;
  assign bpu_io_status_spie = csr_io_status_spie;
  assign bpu_io_status_upie = csr_io_status_upie;
  assign bpu_io_status_mie = csr_io_status_mie;
  assign bpu_io_status_hie = csr_io_status_hie;
  assign bpu_io_status_sie = csr_io_status_sie;
  assign bpu_io_status_uie = csr_io_status_uie;
  assign bpu_io_bp_0_control_ttype = csr_io_bp_0_control_ttype;
  assign bpu_io_bp_0_control_dmode = csr_io_bp_0_control_dmode;
  assign bpu_io_bp_0_control_maskmax = csr_io_bp_0_control_maskmax;
  assign bpu_io_bp_0_control_reserved = csr_io_bp_0_control_reserved;
  assign bpu_io_bp_0_control_action = csr_io_bp_0_control_action;
  assign bpu_io_bp_0_control_chain = csr_io_bp_0_control_chain;
  assign bpu_io_bp_0_control_zero = csr_io_bp_0_control_zero;
  assign bpu_io_bp_0_control_tmatch = csr_io_bp_0_control_tmatch;
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m;
  assign bpu_io_bp_0_control_h = csr_io_bp_0_control_h;
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s;
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u;
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x;
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w;
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r;
  assign bpu_io_bp_0_address = csr_io_bp_0_address;
  assign bpu_io_pc = ibuf_io_pc[38:0];
  assign bpu_io_ea = mem_reg_wdata[38:0];
  assign id_xcpt_if = ibuf_io_inst_0_bits_pf0 | ibuf_io_inst_0_bits_pf1;
  assign T_7402 = csr_io_interrupt | bpu_io_debug_if;
  assign T_7403 = T_7402 | bpu_io_xcpt_if;
  assign T_7404 = T_7403 | id_xcpt_if;
  assign id_xcpt = T_7404 | id_illegal_insn;
  assign T_7405 = id_xcpt_if ? 2'h1 : 2'h2;
  assign T_7406 = bpu_io_xcpt_if ? 2'h3 : T_7405;
  assign T_7407 = bpu_io_debug_if ? 4'hd : {{2'd0}, T_7406};
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : {{60'd0}, T_7407};
  assign ex_waddr = ex_reg_inst[11:7];
  assign mem_waddr = mem_reg_inst[11:7];
  assign wb_waddr = wb_reg_inst[11:7];
  assign T_7411 = ex_reg_valid & ex_ctrl_wxd;
  assign T_7412 = mem_reg_valid & mem_ctrl_wxd;
  assign T_7414 = mem_ctrl_mem == 1'h0;
  assign T_7415 = T_7412 & T_7414;
  assign T_7417 = 5'h0 == ibuf_io_inst_0_bits_inst_rs1;
  assign T_7418 = ex_waddr == ibuf_io_inst_0_bits_inst_rs1;
  assign id_bypass_src_0_1 = T_7411 & T_7418;
  assign T_7419 = mem_waddr == ibuf_io_inst_0_bits_inst_rs1;
  assign id_bypass_src_0_2 = T_7415 & T_7419;
  assign id_bypass_src_0_3 = T_7412 & T_7419;
  assign T_7421 = 5'h0 == ibuf_io_inst_0_bits_inst_rs2;
  assign T_7422 = ex_waddr == ibuf_io_inst_0_bits_inst_rs2;
  assign id_bypass_src_1_1 = T_7411 & T_7422;
  assign T_7423 = mem_waddr == ibuf_io_inst_0_bits_inst_rs2;
  assign id_bypass_src_1_2 = T_7415 & T_7423;
  assign id_bypass_src_1_3 = T_7412 & T_7423;
  assign bypass_mux_0 = 64'h0;
  assign bypass_mux_1 = mem_reg_wdata;
  assign bypass_mux_2 = wb_reg_wdata;
  assign bypass_mux_3 = io_dmem_resp_bits_data_word_bypass;
  assign T_7452 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0};
  assign GEN_0 = GEN_4;
  assign GEN_2 = 2'h1 == ex_reg_rs_lsb_0 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_3 = 2'h2 == ex_reg_rs_lsb_0 ? bypass_mux_2 : GEN_2;
  assign GEN_4 = 2'h3 == ex_reg_rs_lsb_0 ? bypass_mux_3 : GEN_3;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? GEN_0 : T_7452;
  assign T_7453 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1};
  assign GEN_1 = GEN_7;
  assign GEN_5 = 2'h1 == ex_reg_rs_lsb_1 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_6 = 2'h2 == ex_reg_rs_lsb_1 ? bypass_mux_2 : GEN_5;
  assign GEN_7 = 2'h3 == ex_reg_rs_lsb_1 ? bypass_mux_3 : GEN_6;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? GEN_1 : T_7453;
  assign T_7454 = ex_ctrl_sel_imm == 3'h5;
  assign T_7456 = ex_reg_inst[31];
  assign T_7457 = $signed(T_7456);
  assign T_7458 = T_7454 ? $signed(1'sh0) : $signed(T_7457);
  assign T_7459 = ex_ctrl_sel_imm == 3'h2;
  assign T_7460 = ex_reg_inst[30:20];
  assign T_7461 = $signed(T_7460);
  assign T_7462 = T_7459 ? $signed(T_7461) : $signed({11{T_7458}});
  assign T_7463 = ex_ctrl_sel_imm != 3'h2;
  assign T_7464 = ex_ctrl_sel_imm != 3'h3;
  assign T_7465 = T_7463 & T_7464;
  assign T_7466 = ex_reg_inst[19:12];
  assign T_7467 = $signed(T_7466);
  assign T_7468 = T_7465 ? $signed({8{T_7458}}) : $signed(T_7467);
  assign T_7471 = T_7459 | T_7454;
  assign T_7473 = ex_ctrl_sel_imm == 3'h3;
  assign T_7474 = ex_reg_inst[20];
  assign T_7475 = $signed(T_7474);
  assign T_7476 = ex_ctrl_sel_imm == 3'h1;
  assign T_7477 = ex_reg_inst[7];
  assign T_7478 = $signed(T_7477);
  assign T_7479 = T_7476 ? $signed(T_7478) : $signed(T_7458);
  assign T_7480 = T_7473 ? $signed(T_7475) : $signed(T_7479);
  assign T_7481 = T_7471 ? $signed(1'sh0) : $signed(T_7480);
  assign T_7486 = ex_reg_inst[30:25];
  assign T_7487 = T_7471 ? 6'h0 : T_7486;
  assign T_7490 = ex_ctrl_sel_imm == 3'h0;
  assign T_7492 = T_7490 | T_7476;
  assign T_7493 = ex_reg_inst[11:8];
  assign T_7495 = ex_reg_inst[19:16];
  assign T_7496 = ex_reg_inst[24:21];
  assign T_7497 = T_7454 ? T_7495 : T_7496;
  assign T_7498 = T_7492 ? T_7493 : T_7497;
  assign T_7499 = T_7459 ? 4'h0 : T_7498;
  assign T_7502 = ex_ctrl_sel_imm == 3'h4;
  assign T_7505 = ex_reg_inst[15];
  assign T_7508 = T_7454 ? T_7505 : 1'h0;
  assign T_7510 = T_7502 ? T_7474 : T_7508;
  assign T_7512 = T_7490 ? T_7477 : T_7510;
  assign T_7513 = {T_7487,T_7499};
  assign T_7514 = {T_7513,T_7512};
  assign T_7515 = $unsigned(T_7481);
  assign T_7516 = $unsigned(T_7468);
  assign T_7517 = {T_7516,T_7515};
  assign T_7518 = $unsigned(T_7462);
  assign T_7519 = $unsigned(T_7458);
  assign T_7520 = {T_7519,T_7518};
  assign T_7521 = {T_7520,T_7517};
  assign T_7522 = {T_7521,T_7514};
  assign ex_imm = $signed(T_7522);
  assign T_7524 = $signed(ex_rs_0);
  assign T_7525 = $signed(ex_reg_pc);
  assign T_7526 = 2'h2 == ex_ctrl_sel_alu1;
  assign T_7527 = T_7526 ? $signed(T_7525) : $signed(40'sh0);
  assign T_7528 = 2'h1 == ex_ctrl_sel_alu1;
  assign ex_op1 = T_7528 ? $signed(T_7524) : $signed({{24{T_7527[39]}},T_7527});
  assign T_7530 = $signed(ex_rs_1);
  assign T_7533 = ex_reg_rvc ? $signed(4'sh2) : $signed(4'sh4);
  assign T_7534 = 2'h1 == ex_ctrl_sel_alu2;
  assign T_7535 = T_7534 ? $signed(T_7533) : $signed(4'sh0);
  assign T_7536 = 2'h3 == ex_ctrl_sel_alu2;
  assign T_7537 = T_7536 ? $signed(ex_imm) : $signed({{28{T_7535[3]}},T_7535});
  assign T_7538 = 2'h2 == ex_ctrl_sel_alu2;
  assign ex_op2 = T_7538 ? $signed(T_7530) : $signed({{32{T_7537[31]}},T_7537});
  assign alu_clk = clk;
  assign alu_reset = reset;
  assign alu_io_dw = ex_ctrl_alu_dw;
  assign alu_io_fn = ex_ctrl_alu_fn;
  assign alu_io_in2 = T_7539;
  assign alu_io_in1 = T_7540;
  assign T_7539 = $unsigned(ex_op2);
  assign T_7540 = $unsigned(ex_op1);
  assign div_clk = clk;
  assign div_reset = reset;
  assign div_io_req_valid = T_7541;
  assign div_io_req_bits_fn = ex_ctrl_alu_fn;
  assign div_io_req_bits_dw = ex_ctrl_alu_dw;
  assign div_io_req_bits_in1 = ex_rs_0;
  assign div_io_req_bits_in2 = ex_rs_1;
  assign div_io_req_bits_tag = ex_waddr;
  assign div_io_kill = T_7897;
  assign div_io_resp_ready = GEN_150;
  assign T_7541 = ex_reg_valid & ex_ctrl_div;
  assign T_7543 = ctrl_killd == 1'h0;
  assign T_7545 = take_pc_mem_wb == 1'h0;
  assign T_7546 = T_7545 & ibuf_io_inst_0_valid;
  assign T_7547 = T_7546 & ibuf_io_inst_0_bits_replay;
  assign T_7550 = T_7543 & id_xcpt;
  assign T_7554 = T_7546 & csr_io_interrupt;
  assign GEN_8 = id_xcpt ? id_cause : ex_reg_cause;
  assign GEN_9 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_taken : ex_reg_btb_resp_taken;
  assign GEN_10 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_mask : ex_reg_btb_resp_mask;
  assign GEN_11 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_bridx : ex_reg_btb_resp_bridx;
  assign GEN_12 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_target : ex_reg_btb_resp_target;
  assign GEN_13 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_entry : ex_reg_btb_resp_entry;
  assign GEN_14 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_bht_history : ex_reg_btb_resp_bht_history;
  assign GEN_15 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_bht_value : ex_reg_btb_resp_bht_value;
  assign T_7558 = bpu_io_xcpt_if == 1'h0;
  assign T_7560 = ibuf_io_inst_0_bits_pf0 == 1'h0;
  assign T_7561 = T_7558 & T_7560;
  assign T_7562 = T_7561 & ibuf_io_inst_0_bits_pf1;
  assign GEN_16 = T_7562 ? 2'h1 : 2'h0;
  assign GEN_17 = T_7562 ? 1'h1 : ibuf_io_inst_0_bits_rvc;
  assign GEN_18 = id_xcpt ? 4'h0 : id_ctrl_alu_fn;
  assign GEN_19 = id_xcpt ? 1'h1 : id_ctrl_alu_dw;
  assign GEN_20 = id_xcpt ? 2'h2 : id_ctrl_sel_alu1;
  assign GEN_21 = id_xcpt ? GEN_16 : id_ctrl_sel_alu2;
  assign GEN_22 = id_xcpt ? GEN_17 : ibuf_io_inst_0_bits_rvc;
  assign T_7564 = id_ctrl_fence_i | id_csr_flush;
  assign T_7565 = T_7564 | csr_io_singleStep;
  assign T_7566 = id_ctrl_jalr & csr_io_status_debug;
  assign GEN_23 = T_7566 ? 1'h1 : T_7565;
  assign GEN_24 = T_7566 ? 1'h1 : id_ctrl_fence_i;
  assign T_7569 = T_7417 | id_bypass_src_0_1;
  assign T_7570 = T_7569 | id_bypass_src_0_2;
  assign T_7571 = T_7570 | id_bypass_src_0_3;
  assign T_7576 = id_bypass_src_0_2 ? 2'h2 : 2'h3;
  assign T_7577 = id_bypass_src_0_1 ? 2'h1 : T_7576;
  assign T_7578 = T_7417 ? 2'h0 : T_7577;
  assign T_7580 = T_7571 == 1'h0;
  assign T_7581 = id_ctrl_rxs1 & T_7580;
  assign T_7582 = id_rs_0[1:0];
  assign T_7583 = id_rs_0[63:2];
  assign GEN_25 = T_7581 ? T_7582 : T_7578;
  assign GEN_26 = T_7581 ? T_7583 : ex_reg_rs_msb_0;
  assign T_7584 = T_7421 | id_bypass_src_1_1;
  assign T_7585 = T_7584 | id_bypass_src_1_2;
  assign T_7586 = T_7585 | id_bypass_src_1_3;
  assign T_7591 = id_bypass_src_1_2 ? 2'h2 : 2'h3;
  assign T_7592 = id_bypass_src_1_1 ? 2'h1 : T_7591;
  assign T_7593 = T_7421 ? 2'h0 : T_7592;
  assign T_7595 = T_7586 == 1'h0;
  assign T_7596 = id_ctrl_rxs2 & T_7595;
  assign T_7597 = id_rs_1[1:0];
  assign T_7598 = id_rs_1[63:2];
  assign GEN_27 = T_7596 ? T_7597 : T_7593;
  assign GEN_28 = T_7596 ? T_7598 : ex_reg_rs_msb_1;
  assign GEN_29 = T_7543 ? id_ctrl_legal : ex_ctrl_legal;
  assign GEN_30 = T_7543 ? id_ctrl_fp : ex_ctrl_fp;
  assign GEN_31 = T_7543 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign GEN_32 = T_7543 ? id_ctrl_branch : ex_ctrl_branch;
  assign GEN_33 = T_7543 ? id_ctrl_jal : ex_ctrl_jal;
  assign GEN_34 = T_7543 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign GEN_35 = T_7543 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign GEN_36 = T_7543 ? id_ctrl_rxs1 : ex_ctrl_rxs1;
  assign GEN_37 = T_7543 ? GEN_21 : ex_ctrl_sel_alu2;
  assign GEN_38 = T_7543 ? GEN_20 : ex_ctrl_sel_alu1;
  assign GEN_39 = T_7543 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign GEN_40 = T_7543 ? GEN_19 : ex_ctrl_alu_dw;
  assign GEN_41 = T_7543 ? GEN_18 : ex_ctrl_alu_fn;
  assign GEN_42 = T_7543 ? id_ctrl_mem : ex_ctrl_mem;
  assign GEN_43 = T_7543 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign GEN_44 = T_7543 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign GEN_45 = T_7543 ? id_ctrl_rfs1 : ex_ctrl_rfs1;
  assign GEN_46 = T_7543 ? id_ctrl_rfs2 : ex_ctrl_rfs2;
  assign GEN_47 = T_7543 ? id_ctrl_rfs3 : ex_ctrl_rfs3;
  assign GEN_48 = T_7543 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign GEN_49 = T_7543 ? id_ctrl_div : ex_ctrl_div;
  assign GEN_50 = T_7543 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign GEN_51 = T_7543 ? id_csr : ex_ctrl_csr;
  assign GEN_52 = T_7543 ? GEN_24 : ex_ctrl_fence_i;
  assign GEN_53 = T_7543 ? id_ctrl_fence : ex_ctrl_fence;
  assign GEN_54 = T_7543 ? id_ctrl_amo : ex_ctrl_amo;
  assign GEN_55 = T_7543 ? GEN_22 : ex_reg_rvc;
  assign GEN_56 = T_7543 ? GEN_23 : ex_reg_flush_pipe;
  assign GEN_57 = T_7543 ? id_load_use : ex_reg_load_use;
  assign GEN_58 = T_7543 ? T_7571 : ex_reg_rs_bypass_0;
  assign GEN_59 = T_7543 ? GEN_25 : ex_reg_rs_lsb_0;
  assign GEN_60 = T_7543 ? GEN_26 : ex_reg_rs_msb_0;
  assign GEN_61 = T_7543 ? T_7586 : ex_reg_rs_bypass_1;
  assign GEN_62 = T_7543 ? GEN_27 : ex_reg_rs_lsb_1;
  assign GEN_63 = T_7543 ? GEN_28 : ex_reg_rs_msb_1;
  assign T_7601 = T_7543 | csr_io_interrupt;
  assign T_7602 = T_7601 | ibuf_io_inst_0_bits_replay;
  assign GEN_64 = T_7602 ? ibuf_io_inst_0_bits_inst_bits : ex_reg_inst;
  assign GEN_65 = T_7602 ? ibuf_io_pc : ex_reg_pc;
  assign T_7603 = ex_reg_valid | ex_reg_replay;
  assign ex_pc_valid = T_7603 | ex_reg_xcpt_interrupt;
  assign T_7605 = io_dmem_resp_valid == 1'h0;
  assign wb_dcache_miss = wb_ctrl_mem & T_7605;
  assign T_7607 = io_dmem_req_ready == 1'h0;
  assign T_7608 = ex_ctrl_mem & T_7607;
  assign T_7610 = div_io_req_ready == 1'h0;
  assign T_7611 = ex_ctrl_div & T_7610;
  assign replay_ex_structural = T_7608 | T_7611;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T_7612 = replay_ex_structural | replay_ex_load_use;
  assign T_7613 = ex_reg_valid & T_7612;
  assign replay_ex = ex_reg_replay | T_7613;
  assign T_7614 = take_pc_mem_wb | replay_ex;
  assign T_7616 = ex_reg_valid == 1'h0;
  assign ctrl_killx = T_7614 | T_7616;
  assign T_7617 = ex_ctrl_mem_cmd == 5'h7;
  assign T_7623_0 = 3'h0;
  assign T_7623_1 = 3'h4;
  assign T_7623_2 = 3'h1;
  assign T_7623_3 = 3'h5;
  assign T_7625 = T_7623_0 == ex_ctrl_mem_type;
  assign T_7626 = T_7623_1 == ex_ctrl_mem_type;
  assign T_7627 = T_7623_2 == ex_ctrl_mem_type;
  assign T_7628 = T_7623_3 == ex_ctrl_mem_type;
  assign T_7631 = T_7625 | T_7626;
  assign T_7632 = T_7631 | T_7627;
  assign T_7633 = T_7632 | T_7628;
  assign ex_slow_bypass = T_7617 | T_7633;
  assign T_7634 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T_7635 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign ex_xcpt = T_7634 | T_7635;
  assign ex_cause = T_7634 ? ex_reg_cause : 64'h2;
  assign mem_br_taken = mem_reg_wdata[0];
  assign T_7637 = $signed(mem_reg_pc);
  assign T_7638 = mem_ctrl_branch & mem_br_taken;
  assign T_7641 = mem_reg_inst[31];
  assign T_7642 = $signed(T_7641);
  assign T_7647 = {11{T_7642}};
  assign T_7651 = mem_reg_inst[19:12];
  assign T_7652 = $signed(T_7651);
  assign T_7653 = {8{T_7642}};
  assign T_7659 = mem_reg_inst[20];
  assign T_7660 = $signed(T_7659);
  assign T_7662 = mem_reg_inst[7];
  assign T_7663 = $signed(T_7662);
  assign T_7671 = mem_reg_inst[30:25];
  assign T_7678 = mem_reg_inst[11:8];
  assign T_7681 = mem_reg_inst[24:21];
  assign T_7698 = {T_7671,T_7678};
  assign T_7699 = {T_7698,1'h0};
  assign T_7700 = $unsigned(T_7663);
  assign T_7701 = $unsigned(T_7653);
  assign T_7702 = {T_7701,T_7700};
  assign T_7703 = $unsigned(T_7647);
  assign T_7704 = $unsigned(T_7642);
  assign T_7705 = {T_7704,T_7703};
  assign T_7706 = {T_7705,T_7702};
  assign T_7707 = {T_7706,T_7699};
  assign T_7708 = $signed(T_7707);
  assign T_7768 = {T_7671,T_7681};
  assign T_7769 = {T_7768,1'h0};
  assign T_7770 = $unsigned(T_7660);
  assign T_7771 = $unsigned(T_7652);
  assign T_7772 = {T_7771,T_7770};
  assign T_7776 = {T_7705,T_7772};
  assign T_7777 = {T_7776,T_7769};
  assign T_7778 = $signed(T_7777);
  assign T_7781 = mem_reg_rvc ? $signed(4'sh2) : $signed(4'sh4);
  assign T_7782 = mem_ctrl_jal ? $signed(T_7778) : $signed({{28{T_7781[3]}},T_7781});
  assign T_7783 = T_7638 ? $signed(T_7708) : $signed(T_7782);
  assign GEN_171 = {{8{T_7783[31]}},T_7783};
  assign T_7784 = $signed(T_7637) + $signed(GEN_171);
  assign T_7785 = T_7784[39:0];
  assign mem_br_target = $signed(T_7785);
  assign T_7786 = mem_reg_wdata[63:38];
  assign T_7787 = mem_reg_wdata[39:38];
  assign T_7788 = $signed(T_7787);
  assign T_7790 = T_7786 == 26'h0;
  assign T_7792 = T_7786 == 26'h1;
  assign T_7793 = T_7790 | T_7792;
  assign T_7795 = $signed(T_7788) != $signed(2'sh0);
  assign T_7796 = $signed(T_7786);
  assign T_7798 = $signed(T_7796) == $signed(26'sh3ffffff);
  assign T_7801 = $signed(T_7796) == $signed(26'sh3fffffe);
  assign T_7802 = T_7798 | T_7801;
  assign T_7804 = $signed(T_7788) == $signed(2'sh3);
  assign T_7805 = T_7788[0];
  assign T_7806 = T_7802 ? T_7804 : T_7805;
  assign T_7807 = T_7793 ? T_7795 : T_7806;
  assign T_7808 = mem_reg_wdata[38:0];
  assign T_7809 = {T_7807,T_7808};
  assign T_7810 = $signed(T_7809);
  assign T_7811 = mem_ctrl_jalr ? $signed(T_7810) : $signed(mem_br_target);
  assign T_7813 = $signed(T_7811) & $signed(40'shfffffffffe);
  assign T_7814 = $signed(T_7813);
  assign mem_npc = $unsigned(T_7814);
  assign T_7815 = mem_npc != ex_reg_pc;
  assign T_7816 = mem_npc != ibuf_io_pc;
  assign T_7818 = ibuf_io_inst_0_valid ? T_7816 : 1'h1;
  assign mem_wrong_npc = ex_pc_valid ? T_7815 : T_7818;
  assign T_7820 = mem_reg_xcpt == 1'h0;
  assign T_7822 = T_7820 & mem_ctrl_jalr;
  assign T_7823 = $signed(mem_reg_wdata);
  assign T_7824 = T_7822 ? $signed({{24{mem_br_target[39]}},mem_br_target}) : $signed(T_7823);
  assign mem_int_wdata = $unsigned(T_7824);
  assign T_7825 = mem_ctrl_branch | mem_ctrl_jalr;
  assign mem_cfi = T_7825 | mem_ctrl_jal;
  assign T_7827 = T_7638 | mem_ctrl_jalr;
  assign mem_misprediction = T_7827 | mem_ctrl_jal;
  assign T_7828 = mem_misprediction | mem_reg_flush_pipe;
  assign T_7829 = mem_reg_valid & T_7828;
  assign T_7831 = ctrl_killx == 1'h0;
  assign T_7834 = T_7545 & replay_ex;
  assign T_7837 = T_7831 & ex_xcpt;
  assign T_7840 = T_7545 & ex_reg_xcpt_interrupt;
  assign GEN_66 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign T_7841 = ex_ctrl_mem_cmd == 5'h0;
  assign T_7842 = ex_ctrl_mem_cmd == 5'h6;
  assign T_7843 = T_7841 | T_7842;
  assign T_7845 = T_7843 | T_7617;
  assign T_7846 = ex_ctrl_mem_cmd[3];
  assign T_7847 = ex_ctrl_mem_cmd == 5'h4;
  assign T_7848 = T_7846 | T_7847;
  assign T_7849 = T_7845 | T_7848;
  assign T_7850 = ex_ctrl_mem & T_7849;
  assign T_7851 = ex_ctrl_mem_cmd == 5'h1;
  assign T_7853 = T_7851 | T_7617;
  assign T_7857 = T_7853 | T_7848;
  assign T_7858 = ex_ctrl_mem & T_7857;
  assign GEN_67 = ex_reg_btb_hit ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign GEN_68 = ex_reg_btb_hit ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign GEN_69 = ex_reg_btb_hit ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign GEN_70 = ex_reg_btb_hit ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign GEN_71 = ex_reg_btb_hit ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign GEN_72 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign GEN_73 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T_7859 = ex_ctrl_mem | ex_ctrl_rocc;
  assign T_7860 = ex_ctrl_rxs2 & T_7859;
  assign GEN_74 = T_7860 ? ex_rs_1 : mem_reg_rs2;
  assign GEN_75 = ex_pc_valid ? ex_ctrl_legal : mem_ctrl_legal;
  assign GEN_76 = ex_pc_valid ? ex_ctrl_fp : mem_ctrl_fp;
  assign GEN_77 = ex_pc_valid ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign GEN_78 = ex_pc_valid ? ex_ctrl_branch : mem_ctrl_branch;
  assign GEN_79 = ex_pc_valid ? ex_ctrl_jal : mem_ctrl_jal;
  assign GEN_80 = ex_pc_valid ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign GEN_81 = ex_pc_valid ? ex_ctrl_rxs2 : mem_ctrl_rxs2;
  assign GEN_82 = ex_pc_valid ? ex_ctrl_rxs1 : mem_ctrl_rxs1;
  assign GEN_83 = ex_pc_valid ? ex_ctrl_sel_alu2 : mem_ctrl_sel_alu2;
  assign GEN_84 = ex_pc_valid ? ex_ctrl_sel_alu1 : mem_ctrl_sel_alu1;
  assign GEN_85 = ex_pc_valid ? ex_ctrl_sel_imm : mem_ctrl_sel_imm;
  assign GEN_86 = ex_pc_valid ? ex_ctrl_alu_dw : mem_ctrl_alu_dw;
  assign GEN_87 = ex_pc_valid ? ex_ctrl_alu_fn : mem_ctrl_alu_fn;
  assign GEN_88 = ex_pc_valid ? ex_ctrl_mem : mem_ctrl_mem;
  assign GEN_89 = ex_pc_valid ? ex_ctrl_mem_cmd : mem_ctrl_mem_cmd;
  assign GEN_90 = ex_pc_valid ? ex_ctrl_mem_type : mem_ctrl_mem_type;
  assign GEN_91 = ex_pc_valid ? ex_ctrl_rfs1 : mem_ctrl_rfs1;
  assign GEN_92 = ex_pc_valid ? ex_ctrl_rfs2 : mem_ctrl_rfs2;
  assign GEN_93 = ex_pc_valid ? ex_ctrl_rfs3 : mem_ctrl_rfs3;
  assign GEN_94 = ex_pc_valid ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign GEN_95 = ex_pc_valid ? ex_ctrl_div : mem_ctrl_div;
  assign GEN_96 = ex_pc_valid ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign GEN_97 = ex_pc_valid ? ex_ctrl_csr : mem_ctrl_csr;
  assign GEN_98 = ex_pc_valid ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign GEN_99 = ex_pc_valid ? ex_ctrl_fence : mem_ctrl_fence;
  assign GEN_100 = ex_pc_valid ? ex_ctrl_amo : mem_ctrl_amo;
  assign GEN_101 = ex_pc_valid ? ex_reg_rvc : mem_reg_rvc;
  assign GEN_102 = ex_pc_valid ? T_7850 : mem_reg_load;
  assign GEN_103 = ex_pc_valid ? T_7858 : mem_reg_store;
  assign GEN_104 = ex_pc_valid ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign GEN_105 = ex_pc_valid ? GEN_67 : mem_reg_btb_resp_taken;
  assign GEN_106 = ex_pc_valid ? GEN_68 : mem_reg_btb_resp_mask;
  assign GEN_107 = ex_pc_valid ? GEN_69 : mem_reg_btb_resp_bridx;
  assign GEN_108 = ex_pc_valid ? GEN_70 : mem_reg_btb_resp_target;
  assign GEN_109 = ex_pc_valid ? GEN_71 : mem_reg_btb_resp_entry;
  assign GEN_110 = ex_pc_valid ? GEN_72 : mem_reg_btb_resp_bht_history;
  assign GEN_111 = ex_pc_valid ? GEN_73 : mem_reg_btb_resp_bht_value;
  assign GEN_112 = ex_pc_valid ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign GEN_113 = ex_pc_valid ? ex_slow_bypass : mem_reg_slow_bypass;
  assign GEN_114 = ex_pc_valid ? ex_reg_inst : mem_reg_inst;
  assign GEN_115 = ex_pc_valid ? ex_reg_pc : mem_reg_pc;
  assign GEN_116 = ex_pc_valid ? alu_io_out : mem_reg_wdata;
  assign GEN_117 = ex_pc_valid ? GEN_74 : mem_reg_rs2;
  assign T_7861 = mem_reg_load & bpu_io_xcpt_ld;
  assign T_7862 = mem_reg_store & bpu_io_xcpt_st;
  assign mem_breakpoint = T_7861 | T_7862;
  assign T_7863 = mem_reg_load & bpu_io_debug_ld;
  assign T_7864 = mem_reg_store & bpu_io_debug_st;
  assign mem_debug_breakpoint = T_7863 | T_7864;
  assign T_7868 = mem_ctrl_mem & io_dmem_xcpt_ma_st;
  assign T_7870 = mem_ctrl_mem & io_dmem_xcpt_ma_ld;
  assign T_7872 = mem_ctrl_mem & io_dmem_xcpt_pf_st;
  assign T_7874 = mem_ctrl_mem & io_dmem_xcpt_pf_ld;
  assign T_7876 = mem_debug_breakpoint | mem_breakpoint;
  assign T_7878 = T_7876 | T_7868;
  assign T_7879 = T_7878 | T_7870;
  assign T_7880 = T_7879 | T_7872;
  assign mem_new_xcpt = T_7880 | T_7874;
  assign T_7881 = T_7872 ? 3'h7 : 3'h5;
  assign T_7882 = T_7870 ? 3'h4 : T_7881;
  assign T_7883 = T_7868 ? 3'h6 : T_7882;
  assign T_7885 = mem_breakpoint ? 3'h3 : T_7883;
  assign mem_new_cause = mem_debug_breakpoint ? 4'hd : {{1'd0}, T_7885};
  assign T_7886 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T_7887 = mem_reg_valid & mem_new_xcpt;
  assign mem_xcpt = T_7886 | T_7887;
  assign mem_cause = T_7886 ? mem_reg_cause : {{60'd0}, mem_new_cause};
  assign dcache_kill_mem = T_7412 & io_dmem_replay_next;
  assign T_7889 = mem_reg_valid & mem_ctrl_fp;
  assign fpu_kill_mem = T_7889 & io_fpu_nack_mem;
  assign T_7890 = dcache_kill_mem | mem_reg_replay;
  assign replay_mem = T_7890 | fpu_kill_mem;
  assign T_7891 = dcache_kill_mem | take_pc_wb;
  assign T_7892 = T_7891 | mem_reg_xcpt;
  assign T_7894 = mem_reg_valid == 1'h0;
  assign killm_common = T_7892 | T_7894;
  assign T_7895 = div_io_req_ready & div_io_req_valid;
  assign T_7897 = killm_common & T_7896;
  assign T_7898 = killm_common | mem_xcpt;
  assign ctrl_killm = T_7898 | fpu_kill_mem;
  assign T_7900 = ctrl_killm == 1'h0;
  assign T_7902 = take_pc_wb == 1'h0;
  assign T_7903 = replay_mem & T_7902;
  assign T_7906 = mem_xcpt & T_7902;
  assign GEN_118 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign T_7907 = mem_reg_valid | mem_reg_replay;
  assign T_7908 = T_7907 | mem_reg_xcpt_interrupt;
  assign T_7911 = T_7820 & mem_ctrl_fp;
  assign T_7912 = T_7911 & mem_ctrl_wxd;
  assign T_7913 = T_7912 ? io_fpu_toint_data : mem_int_wdata;
  assign GEN_119 = mem_ctrl_rocc ? mem_reg_rs2 : wb_reg_rs2;
  assign GEN_120 = T_7908 ? mem_ctrl_legal : wb_ctrl_legal;
  assign GEN_121 = T_7908 ? mem_ctrl_fp : wb_ctrl_fp;
  assign GEN_122 = T_7908 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign GEN_123 = T_7908 ? mem_ctrl_branch : wb_ctrl_branch;
  assign GEN_124 = T_7908 ? mem_ctrl_jal : wb_ctrl_jal;
  assign GEN_125 = T_7908 ? mem_ctrl_jalr : wb_ctrl_jalr;
  assign GEN_126 = T_7908 ? mem_ctrl_rxs2 : wb_ctrl_rxs2;
  assign GEN_127 = T_7908 ? mem_ctrl_rxs1 : wb_ctrl_rxs1;
  assign GEN_128 = T_7908 ? mem_ctrl_sel_alu2 : wb_ctrl_sel_alu2;
  assign GEN_129 = T_7908 ? mem_ctrl_sel_alu1 : wb_ctrl_sel_alu1;
  assign GEN_130 = T_7908 ? mem_ctrl_sel_imm : wb_ctrl_sel_imm;
  assign GEN_131 = T_7908 ? mem_ctrl_alu_dw : wb_ctrl_alu_dw;
  assign GEN_132 = T_7908 ? mem_ctrl_alu_fn : wb_ctrl_alu_fn;
  assign GEN_133 = T_7908 ? mem_ctrl_mem : wb_ctrl_mem;
  assign GEN_134 = T_7908 ? mem_ctrl_mem_cmd : wb_ctrl_mem_cmd;
  assign GEN_135 = T_7908 ? mem_ctrl_mem_type : wb_ctrl_mem_type;
  assign GEN_136 = T_7908 ? mem_ctrl_rfs1 : wb_ctrl_rfs1;
  assign GEN_137 = T_7908 ? mem_ctrl_rfs2 : wb_ctrl_rfs2;
  assign GEN_138 = T_7908 ? mem_ctrl_rfs3 : wb_ctrl_rfs3;
  assign GEN_139 = T_7908 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign GEN_140 = T_7908 ? mem_ctrl_div : wb_ctrl_div;
  assign GEN_141 = T_7908 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign GEN_142 = T_7908 ? mem_ctrl_csr : wb_ctrl_csr;
  assign GEN_143 = T_7908 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign GEN_144 = T_7908 ? mem_ctrl_fence : wb_ctrl_fence;
  assign GEN_145 = T_7908 ? mem_ctrl_amo : wb_ctrl_amo;
  assign GEN_146 = T_7908 ? T_7913 : wb_reg_wdata;
  assign GEN_147 = T_7908 ? GEN_119 : wb_reg_rs2;
  assign GEN_148 = T_7908 ? mem_reg_inst : wb_reg_inst;
  assign GEN_149 = T_7908 ? mem_reg_pc : wb_reg_pc;
  assign T_7914 = wb_ctrl_div | wb_dcache_miss;
  assign wb_set_sboard = T_7914 | wb_ctrl_rocc;
  assign replay_wb_common = io_dmem_s2_nack | wb_reg_replay;
  assign T_7917 = io_rocc_cmd_ready == 1'h0;
  assign replay_wb_rocc = T_7386 & T_7917;
  assign replay_wb = replay_wb_common | replay_wb_rocc;
  assign wb_xcpt = wb_reg_xcpt | csr_io_csr_xcpt;
  assign T_7918 = replay_wb | wb_xcpt;
  assign T_7919 = T_7918 | csr_io_eret;
  assign T_7920 = io_dmem_resp_bits_tag[0];
  assign dmem_resp_xpu = T_7920 == 1'h0;
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[5:1];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay;
  assign T_7924 = wb_reg_valid & wb_ctrl_wxd;
  assign T_7926 = T_7924 == 1'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign ll_waddr = GEN_151;
  assign T_7927 = div_io_resp_ready & div_io_resp_valid;
  assign ll_wen = GEN_152;
  assign T_7928 = dmem_resp_replay & dmem_resp_xpu;
  assign GEN_150 = T_7928 ? 1'h0 : T_7926;
  assign GEN_151 = T_7928 ? dmem_resp_waddr : div_io_resp_bits_tag;
  assign GEN_152 = T_7928 ? 1'h1 : T_7927;
  assign T_7932 = replay_wb == 1'h0;
  assign T_7933 = wb_reg_valid & T_7932;
  assign T_7935 = wb_xcpt == 1'h0;
  assign wb_valid = T_7933 & T_7935;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign rf_wen = wb_wen | ll_wen;
  assign rf_waddr = ll_wen ? ll_waddr : wb_waddr;
  assign T_7936 = dmem_resp_valid & dmem_resp_xpu;
  assign T_7937 = wb_ctrl_csr != 3'h0;
  assign T_7938 = T_7937 ? csr_io_rw_rdata : wb_reg_wdata;
  assign T_7939 = ll_wen ? ll_wdata : T_7938;
  assign rf_wdata = T_7936 ? io_dmem_resp_bits_data : T_7939;
  assign T_7941 = rf_waddr != 5'h0;
  assign T_7943 = ~ rf_waddr;
  assign T_7945 = rf_waddr == ibuf_io_inst_0_bits_inst_rs1;
  assign GEN_153 = T_7945 ? rf_wdata : T_7202;
  assign T_7946 = rf_waddr == ibuf_io_inst_0_bits_inst_rs2;
  assign GEN_154 = T_7946 ? rf_wdata : T_7212;
  assign GEN_160 = T_7941 ? GEN_153 : T_7202;
  assign GEN_161 = T_7941 ? GEN_154 : T_7212;
  assign GEN_164 = rf_wen ? T_7941 : 1'h0;
  assign GEN_167 = rf_wen ? GEN_160 : T_7202;
  assign GEN_168 = rf_wen ? GEN_161 : T_7212;
  assign T_7947 = wb_reg_wdata[63:38];
  assign T_7948 = wb_reg_wdata[39:38];
  assign T_7949 = $signed(T_7948);
  assign T_7951 = T_7947 == 26'h0;
  assign T_7953 = T_7947 == 26'h1;
  assign T_7954 = T_7951 | T_7953;
  assign T_7956 = $signed(T_7949) != $signed(2'sh0);
  assign T_7957 = $signed(T_7947);
  assign T_7959 = $signed(T_7957) == $signed(26'sh3ffffff);
  assign T_7962 = $signed(T_7957) == $signed(26'sh3fffffe);
  assign T_7963 = T_7959 | T_7962;
  assign T_7965 = $signed(T_7949) == $signed(2'sh3);
  assign T_7966 = T_7949[0];
  assign T_7967 = T_7963 ? T_7965 : T_7966;
  assign T_7968 = T_7954 ? T_7956 : T_7967;
  assign T_7969 = wb_reg_wdata[38:0];
  assign T_7970 = {T_7968,T_7969};
  assign T_7971 = wb_reg_inst[31:20];
  assign T_7972 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign T_7974 = ibuf_io_inst_0_bits_inst_rs1 != 5'h0;
  assign T_7975 = id_ctrl_rxs1 & T_7974;
  assign T_7977 = ibuf_io_inst_0_bits_inst_rs2 != 5'h0;
  assign T_7978 = id_ctrl_rxs2 & T_7977;
  assign T_7980 = ibuf_io_inst_0_bits_inst_rd != 5'h0;
  assign T_7981 = id_ctrl_wxd & T_7980;
  assign T_7984 = T_7983[31:1];
  assign GEN_172 = {{1'd0}, T_7984};
  assign T_7985 = GEN_172 << 1;
  assign T_7988 = 32'h1 << ll_waddr;
  assign T_7990 = ll_wen ? T_7988 : 32'h0;
  assign T_7991 = ~ T_7990;
  assign T_7992 = T_7985 & T_7991;
  assign GEN_169 = ll_wen ? T_7992 : T_7983;
  assign T_7994 = T_7985 >> ibuf_io_inst_0_bits_inst_rs1;
  assign T_7995 = T_7994[0];
  assign T_7996 = T_7975 & T_7995;
  assign T_7997 = T_7985 >> ibuf_io_inst_0_bits_inst_rs2;
  assign T_7998 = T_7997[0];
  assign T_7999 = T_7978 & T_7998;
  assign T_8000 = T_7985 >> ibuf_io_inst_0_bits_inst_rd;
  assign T_8001 = T_8000[0];
  assign T_8002 = T_7981 & T_8001;
  assign T_8003 = T_7996 | T_7999;
  assign id_sboard_hazard = T_8003 | T_8002;
  assign T_8004 = wb_set_sboard & wb_wen;
  assign T_8006 = 32'h1 << wb_waddr;
  assign T_8008 = T_8004 ? T_8006 : 32'h0;
  assign T_8009 = T_7992 | T_8008;
  assign T_8010 = ll_wen | T_8004;
  assign GEN_170 = T_8010 ? T_8009 : GEN_169;
  assign T_8011 = ex_ctrl_csr != 3'h0;
  assign T_8012 = T_8011 | ex_ctrl_jalr;
  assign T_8013 = T_8012 | ex_ctrl_mem;
  assign T_8014 = T_8013 | ex_ctrl_div;
  assign T_8015 = T_8014 | ex_ctrl_fp;
  assign ex_cannot_bypass = T_8015 | ex_ctrl_rocc;
  assign T_8016 = ibuf_io_inst_0_bits_inst_rs1 == ex_waddr;
  assign T_8017 = T_7975 & T_8016;
  assign T_8018 = ibuf_io_inst_0_bits_inst_rs2 == ex_waddr;
  assign T_8019 = T_7978 & T_8018;
  assign T_8020 = ibuf_io_inst_0_bits_inst_rd == ex_waddr;
  assign T_8021 = T_7981 & T_8020;
  assign T_8022 = T_8017 | T_8019;
  assign T_8023 = T_8022 | T_8021;
  assign data_hazard_ex = ex_ctrl_wxd & T_8023;
  assign T_8025 = io_fpu_dec_ren1 & T_8016;
  assign T_8027 = io_fpu_dec_ren2 & T_8018;
  assign T_8028 = ibuf_io_inst_0_bits_inst_rs3 == ex_waddr;
  assign T_8029 = io_fpu_dec_ren3 & T_8028;
  assign T_8031 = io_fpu_dec_wen & T_8020;
  assign T_8032 = T_8025 | T_8027;
  assign T_8033 = T_8032 | T_8029;
  assign T_8034 = T_8033 | T_8031;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T_8034;
  assign T_8035 = data_hazard_ex & ex_cannot_bypass;
  assign T_8036 = T_8035 | fp_data_hazard_ex;
  assign id_ex_hazard = ex_reg_valid & T_8036;
  assign T_8038 = mem_ctrl_csr != 3'h0;
  assign T_8039 = mem_ctrl_mem & mem_reg_slow_bypass;
  assign T_8040 = T_8038 | T_8039;
  assign T_8041 = T_8040 | mem_ctrl_div;
  assign T_8042 = T_8041 | mem_ctrl_fp;
  assign mem_cannot_bypass = T_8042 | mem_ctrl_rocc;
  assign T_8043 = ibuf_io_inst_0_bits_inst_rs1 == mem_waddr;
  assign T_8044 = T_7975 & T_8043;
  assign T_8045 = ibuf_io_inst_0_bits_inst_rs2 == mem_waddr;
  assign T_8046 = T_7978 & T_8045;
  assign T_8047 = ibuf_io_inst_0_bits_inst_rd == mem_waddr;
  assign T_8048 = T_7981 & T_8047;
  assign T_8049 = T_8044 | T_8046;
  assign T_8050 = T_8049 | T_8048;
  assign data_hazard_mem = mem_ctrl_wxd & T_8050;
  assign T_8052 = io_fpu_dec_ren1 & T_8043;
  assign T_8054 = io_fpu_dec_ren2 & T_8045;
  assign T_8055 = ibuf_io_inst_0_bits_inst_rs3 == mem_waddr;
  assign T_8056 = io_fpu_dec_ren3 & T_8055;
  assign T_8058 = io_fpu_dec_wen & T_8047;
  assign T_8059 = T_8052 | T_8054;
  assign T_8060 = T_8059 | T_8056;
  assign T_8061 = T_8060 | T_8058;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T_8061;
  assign T_8062 = data_hazard_mem & mem_cannot_bypass;
  assign T_8063 = T_8062 | fp_data_hazard_mem;
  assign id_mem_hazard = mem_reg_valid & T_8063;
  assign T_8064 = mem_reg_valid & data_hazard_mem;
  assign T_8065 = T_8064 & mem_ctrl_mem;
  assign T_8066 = ibuf_io_inst_0_bits_inst_rs1 == wb_waddr;
  assign T_8067 = T_7975 & T_8066;
  assign T_8068 = ibuf_io_inst_0_bits_inst_rs2 == wb_waddr;
  assign T_8069 = T_7978 & T_8068;
  assign T_8070 = ibuf_io_inst_0_bits_inst_rd == wb_waddr;
  assign T_8071 = T_7981 & T_8070;
  assign T_8072 = T_8067 | T_8069;
  assign T_8073 = T_8072 | T_8071;
  assign data_hazard_wb = wb_ctrl_wxd & T_8073;
  assign T_8075 = io_fpu_dec_ren1 & T_8066;
  assign T_8077 = io_fpu_dec_ren2 & T_8068;
  assign T_8078 = ibuf_io_inst_0_bits_inst_rs3 == wb_waddr;
  assign T_8079 = io_fpu_dec_ren3 & T_8078;
  assign T_8081 = io_fpu_dec_wen & T_8070;
  assign T_8082 = T_8075 | T_8077;
  assign T_8083 = T_8082 | T_8079;
  assign T_8084 = T_8083 | T_8081;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T_8084;
  assign T_8085 = data_hazard_wb & wb_set_sboard;
  assign T_8086 = T_8085 | fp_data_hazard_wb;
  assign id_wb_hazard = wb_reg_valid & T_8086;
  assign T_8090 = io_dmem_req_valid | dcache_blocked;
  assign T_8091 = T_7607 & T_8090;
  assign T_8094 = wb_reg_xcpt == 1'h0;
  assign T_8097 = T_8094 & T_7917;
  assign T_8098 = io_rocc_cmd_valid | rocc_blocked;
  assign T_8099 = T_8097 & T_8098;
  assign T_8100 = id_ex_hazard | id_mem_hazard;
  assign T_8101 = T_8100 | id_wb_hazard;
  assign T_8102 = T_8101 | id_sboard_hazard;
  assign T_8105 = id_ctrl_mem & dcache_blocked;
  assign T_8106 = T_8102 | T_8105;
  assign T_8107 = id_ctrl_rocc & rocc_blocked;
  assign T_8108 = T_8106 | T_8107;
  assign T_8109 = T_8108 | T_7397;
  assign ctrl_stalld = T_8109 | csr_io_csr_stall;
  assign T_8111 = ibuf_io_inst_0_valid == 1'h0;
  assign T_8112 = T_8111 | ibuf_io_inst_0_bits_replay;
  assign T_8113 = T_8112 | take_pc_mem_wb;
  assign T_8114 = T_8113 | ctrl_stalld;
  assign T_8115 = T_8114 | csr_io_interrupt;
  assign T_8118 = wb_xcpt | csr_io_eret;
  assign T_8119 = replay_wb ? wb_reg_pc : mem_npc;
  assign T_8120 = T_8118 ? csr_io_evec : T_8119;
  assign T_8121 = wb_reg_valid & wb_ctrl_fence_i;
  assign T_8123 = io_dmem_s2_nack == 1'h0;
  assign T_8124 = T_8121 & T_8123;
  assign T_8126 = ctrl_stalld == 1'h0;
  assign T_8127 = T_8126 | csr_io_interrupt;
  assign T_8128 = mem_reg_replay & mem_reg_btb_hit;
  assign T_8131 = mem_reg_valid & T_7902;
  assign T_8133 = mem_cfi == 1'h0;
  assign T_8134 = mem_misprediction | T_8133;
  assign T_8135 = T_8131 & T_8134;
  assign T_8136 = T_8135 & mem_wrong_npc;
  assign T_8137 = T_8128 | T_8136;
  assign T_8139 = mem_reg_replay == 1'h0;
  assign T_8140 = T_8139 & mem_cfi;
  assign T_8141 = mem_ctrl_jal | mem_ctrl_jalr;
  assign T_8142 = mem_reg_inst[19:15];
  assign T_8145 = T_8142 & 5'h19;
  assign T_8146 = 5'h1 == T_8145;
  assign T_8147 = mem_ctrl_jalr & T_8146;
  assign T_8150 = mem_reg_rvc ? 2'h0 : 2'h2;
  assign GEN_173 = {{38'd0}, T_8150};
  assign T_8151 = mem_reg_pc + GEN_173;
  assign T_8152 = T_8151[39:0];
  assign T_8153 = ~ io_imem_btb_update_bits_br_pc;
  assign T_8155 = T_8153 | 39'h3;
  assign T_8156 = ~ T_8155;
  assign T_8160 = T_8131 & mem_ctrl_branch;
  assign T_8164 = mem_waddr[0];
  assign T_8165 = io_imem_btb_update_bits_isJump & T_8164;
  assign T_8168 = T_7543 & id_ctrl_fp;
  assign T_8169 = dmem_resp_valid & T_7920;
  assign T_8170 = ex_reg_valid & ex_ctrl_mem;
  assign ex_dcache_tag = {ex_waddr,ex_ctrl_fp};
  assign T_8172 = ex_rs_0[63:38];
  assign T_8173 = alu_io_adder_out[39:38];
  assign T_8174 = $signed(T_8173);
  assign T_8176 = T_8172 == 26'h0;
  assign T_8178 = T_8172 == 26'h1;
  assign T_8179 = T_8176 | T_8178;
  assign T_8181 = $signed(T_8174) != $signed(2'sh0);
  assign T_8182 = $signed(T_8172);
  assign T_8184 = $signed(T_8182) == $signed(26'sh3ffffff);
  assign T_8187 = $signed(T_8182) == $signed(26'sh3fffffe);
  assign T_8188 = T_8184 | T_8187;
  assign T_8190 = $signed(T_8174) == $signed(2'sh3);
  assign T_8191 = T_8174[0];
  assign T_8192 = T_8188 ? T_8190 : T_8191;
  assign T_8193 = T_8179 ? T_8181 : T_8192;
  assign T_8194 = alu_io_adder_out[38:0];
  assign T_8195 = {T_8193,T_8194};
  assign T_8196 = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign T_8197 = killm_common | mem_breakpoint;
  assign T_8199 = io_dmem_s1_kill == 1'h0;
  assign T_8200 = mem_xcpt & T_8199;
  assign T_8201 = {io_dmem_xcpt_pf_ld,io_dmem_xcpt_pf_st};
  assign T_8202 = {io_dmem_xcpt_ma_ld,io_dmem_xcpt_ma_st};
  assign T_8203 = {T_8202,T_8201};
  assign T_8205 = T_8203 != 4'h0;
  assign T_8206 = T_8205 | reset;
  assign T_8208 = T_8206 == 1'h0;
  assign T_8211 = replay_wb_common == 1'h0;
  assign T_8212 = T_7386 & T_8211;
  assign T_8215 = wb_xcpt & T_7374;
  assign T_8234_funct = T_8252;
  assign T_8234_rs2 = T_8251;
  assign T_8234_rs1 = T_8250;
  assign T_8234_xd = T_8249;
  assign T_8234_xs1 = T_8248;
  assign T_8234_xs2 = T_8247;
  assign T_8234_rd = T_8246;
  assign T_8234_opcode = T_8245;
  assign T_8244 = wb_reg_inst;
  assign T_8245 = T_8244[6:0];
  assign T_8246 = T_8244[11:7];
  assign T_8247 = T_8244[12];
  assign T_8248 = T_8244[13];
  assign T_8249 = T_8244[14];
  assign T_8250 = T_8244[19:15];
  assign T_8251 = T_8244[24:20];
  assign T_8252 = T_8244[31:25];
  assign T_8253 = csr_io_time[31:0];
  assign T_8255 = rf_wen ? rf_waddr : 5'h0;
  assign T_8256 = wb_reg_inst[19:15];
  assign T_8259 = wb_reg_inst[24:20];
  assign T_8263 = reset == 1'h0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_155 = GEN_414[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_156 = GEN_415[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_157 = GEN_416[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_158 = GEN_417[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_159 = GEN_418[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_162 = GEN_419[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_163 = GEN_420[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_165 = GEN_421[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_166 = GEN_422[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_174 = GEN_423[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_175 = GEN_424[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_176 = GEN_425[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_177 = GEN_426[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_178 = GEN_427[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_179 = GEN_428[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_180 = GEN_429[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_181 = GEN_430[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_182 = GEN_431[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_183 = GEN_432[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_184 = GEN_433[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_185 = GEN_434[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_186 = GEN_435[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_187 = GEN_436[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_188 = GEN_437[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_189 = GEN_438[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_190 = GEN_439[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_191 = GEN_440[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_192 = GEN_441[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_193 = GEN_442[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_194 = GEN_443[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_195 = GEN_444[39:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_196 = GEN_445[5:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_197 = GEN_446[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_198 = GEN_447[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_199 = GEN_448[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_200 = GEN_449[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_201 = GEN_450[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_202 = GEN_451[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_203 = GEN_452[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_204 = GEN_453[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_205 = GEN_454[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_206 = GEN_455[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_207 = GEN_456[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_208 = GEN_457[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_209 = GEN_458[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_210 = GEN_459[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_211 = GEN_460[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_212 = GEN_461[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_213 = GEN_462[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_214 = GEN_463[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_215 = GEN_464[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_216 = GEN_465[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_217 = GEN_466[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_218 = GEN_467[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_219 = GEN_468[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_220 = GEN_469[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_221 = GEN_470[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_222 = GEN_471[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_223 = GEN_472[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_224 = GEN_473[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_225 = GEN_474[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_226 = GEN_475[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_227 = GEN_476[39:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_228 = GEN_477[5:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_229 = GEN_478[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_230 = GEN_479[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_231 = GEN_480[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_232 = GEN_481[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_233 = GEN_482[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_234 = GEN_483[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_235 = GEN_484[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_236 = GEN_485[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_237 = GEN_486[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_238 = GEN_487[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_239 = GEN_488[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_240 = GEN_489[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_241 = GEN_490[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_242 = GEN_491[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_243 = GEN_492[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_244 = GEN_493[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_245 = GEN_494[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_246 = GEN_495[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_247 = GEN_496[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_248 = GEN_497[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_249 = GEN_498[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_250 = GEN_499[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_251 = GEN_500[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_252 = GEN_501[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_253 = GEN_502[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_254 = GEN_503[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_255 = GEN_504[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_256 = GEN_505[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_257 = GEN_506[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_258 = GEN_507[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_259 = GEN_508[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_260 = GEN_509[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_261 = GEN_510[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_262 = GEN_511[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_263 = GEN_512[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_264 = GEN_513[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_265 = GEN_514[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_266 = GEN_515[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_267 = GEN_516[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_268 = GEN_517[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_269 = GEN_518[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_270 = {1{$random}};
  ex_ctrl_legal = GEN_270[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_271 = {1{$random}};
  ex_ctrl_fp = GEN_271[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_272 = {1{$random}};
  ex_ctrl_rocc = GEN_272[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_273 = {1{$random}};
  ex_ctrl_branch = GEN_273[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_274 = {1{$random}};
  ex_ctrl_jal = GEN_274[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_275 = {1{$random}};
  ex_ctrl_jalr = GEN_275[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_276 = {1{$random}};
  ex_ctrl_rxs2 = GEN_276[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_277 = {1{$random}};
  ex_ctrl_rxs1 = GEN_277[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_278 = {1{$random}};
  ex_ctrl_sel_alu2 = GEN_278[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_279 = {1{$random}};
  ex_ctrl_sel_alu1 = GEN_279[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_280 = {1{$random}};
  ex_ctrl_sel_imm = GEN_280[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_281 = {1{$random}};
  ex_ctrl_alu_dw = GEN_281[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_282 = {1{$random}};
  ex_ctrl_alu_fn = GEN_282[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_283 = {1{$random}};
  ex_ctrl_mem = GEN_283[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_284 = {1{$random}};
  ex_ctrl_mem_cmd = GEN_284[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_285 = {1{$random}};
  ex_ctrl_mem_type = GEN_285[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_286 = {1{$random}};
  ex_ctrl_rfs1 = GEN_286[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_287 = {1{$random}};
  ex_ctrl_rfs2 = GEN_287[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_288 = {1{$random}};
  ex_ctrl_rfs3 = GEN_288[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_289 = {1{$random}};
  ex_ctrl_wfd = GEN_289[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_290 = {1{$random}};
  ex_ctrl_div = GEN_290[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_291 = {1{$random}};
  ex_ctrl_wxd = GEN_291[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_292 = {1{$random}};
  ex_ctrl_csr = GEN_292[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_293 = {1{$random}};
  ex_ctrl_fence_i = GEN_293[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_294 = {1{$random}};
  ex_ctrl_fence = GEN_294[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_295 = {1{$random}};
  ex_ctrl_amo = GEN_295[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_296 = {1{$random}};
  mem_ctrl_legal = GEN_296[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_297 = {1{$random}};
  mem_ctrl_fp = GEN_297[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_298 = {1{$random}};
  mem_ctrl_rocc = GEN_298[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_299 = {1{$random}};
  mem_ctrl_branch = GEN_299[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_300 = {1{$random}};
  mem_ctrl_jal = GEN_300[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_301 = {1{$random}};
  mem_ctrl_jalr = GEN_301[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_302 = {1{$random}};
  mem_ctrl_rxs2 = GEN_302[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_303 = {1{$random}};
  mem_ctrl_rxs1 = GEN_303[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_304 = {1{$random}};
  mem_ctrl_sel_alu2 = GEN_304[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_305 = {1{$random}};
  mem_ctrl_sel_alu1 = GEN_305[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_306 = {1{$random}};
  mem_ctrl_sel_imm = GEN_306[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_307 = {1{$random}};
  mem_ctrl_alu_dw = GEN_307[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_308 = {1{$random}};
  mem_ctrl_alu_fn = GEN_308[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_309 = {1{$random}};
  mem_ctrl_mem = GEN_309[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_310 = {1{$random}};
  mem_ctrl_mem_cmd = GEN_310[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_311 = {1{$random}};
  mem_ctrl_mem_type = GEN_311[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_312 = {1{$random}};
  mem_ctrl_rfs1 = GEN_312[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_313 = {1{$random}};
  mem_ctrl_rfs2 = GEN_313[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_314 = {1{$random}};
  mem_ctrl_rfs3 = GEN_314[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_315 = {1{$random}};
  mem_ctrl_wfd = GEN_315[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_316 = {1{$random}};
  mem_ctrl_div = GEN_316[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_317 = {1{$random}};
  mem_ctrl_wxd = GEN_317[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_318 = {1{$random}};
  mem_ctrl_csr = GEN_318[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_319 = {1{$random}};
  mem_ctrl_fence_i = GEN_319[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_320 = {1{$random}};
  mem_ctrl_fence = GEN_320[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_321 = {1{$random}};
  mem_ctrl_amo = GEN_321[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_322 = {1{$random}};
  wb_ctrl_legal = GEN_322[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_323 = {1{$random}};
  wb_ctrl_fp = GEN_323[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_324 = {1{$random}};
  wb_ctrl_rocc = GEN_324[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_325 = {1{$random}};
  wb_ctrl_branch = GEN_325[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_326 = {1{$random}};
  wb_ctrl_jal = GEN_326[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_327 = {1{$random}};
  wb_ctrl_jalr = GEN_327[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_328 = {1{$random}};
  wb_ctrl_rxs2 = GEN_328[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_329 = {1{$random}};
  wb_ctrl_rxs1 = GEN_329[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_330 = {1{$random}};
  wb_ctrl_sel_alu2 = GEN_330[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_331 = {1{$random}};
  wb_ctrl_sel_alu1 = GEN_331[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_332 = {1{$random}};
  wb_ctrl_sel_imm = GEN_332[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_333 = {1{$random}};
  wb_ctrl_alu_dw = GEN_333[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_334 = {1{$random}};
  wb_ctrl_alu_fn = GEN_334[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_335 = {1{$random}};
  wb_ctrl_mem = GEN_335[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_336 = {1{$random}};
  wb_ctrl_mem_cmd = GEN_336[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_337 = {1{$random}};
  wb_ctrl_mem_type = GEN_337[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_338 = {1{$random}};
  wb_ctrl_rfs1 = GEN_338[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_339 = {1{$random}};
  wb_ctrl_rfs2 = GEN_339[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_340 = {1{$random}};
  wb_ctrl_rfs3 = GEN_340[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_341 = {1{$random}};
  wb_ctrl_wfd = GEN_341[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_342 = {1{$random}};
  wb_ctrl_div = GEN_342[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_343 = {1{$random}};
  wb_ctrl_wxd = GEN_343[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_344 = {1{$random}};
  wb_ctrl_csr = GEN_344[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_345 = {1{$random}};
  wb_ctrl_fence_i = GEN_345[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_346 = {1{$random}};
  wb_ctrl_fence = GEN_346[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_347 = {1{$random}};
  wb_ctrl_amo = GEN_347[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_348 = {1{$random}};
  ex_reg_xcpt_interrupt = GEN_348[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_349 = {1{$random}};
  ex_reg_valid = GEN_349[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_350 = {1{$random}};
  ex_reg_rvc = GEN_350[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_351 = {1{$random}};
  ex_reg_btb_hit = GEN_351[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_352 = {1{$random}};
  ex_reg_btb_resp_taken = GEN_352[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_353 = {1{$random}};
  ex_reg_btb_resp_mask = GEN_353[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_354 = {1{$random}};
  ex_reg_btb_resp_bridx = GEN_354[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_355 = {2{$random}};
  ex_reg_btb_resp_target = GEN_355[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_356 = {1{$random}};
  ex_reg_btb_resp_entry = GEN_356[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_357 = {1{$random}};
  ex_reg_btb_resp_bht_history = GEN_357[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_358 = {1{$random}};
  ex_reg_btb_resp_bht_value = GEN_358[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_359 = {1{$random}};
  ex_reg_xcpt = GEN_359[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_360 = {1{$random}};
  ex_reg_flush_pipe = GEN_360[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_361 = {1{$random}};
  ex_reg_load_use = GEN_361[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_362 = {2{$random}};
  ex_reg_cause = GEN_362[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_363 = {1{$random}};
  ex_reg_replay = GEN_363[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_364 = {2{$random}};
  ex_reg_pc = GEN_364[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_365 = {1{$random}};
  ex_reg_inst = GEN_365[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_366 = {1{$random}};
  mem_reg_xcpt_interrupt = GEN_366[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_367 = {1{$random}};
  mem_reg_valid = GEN_367[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_368 = {1{$random}};
  mem_reg_rvc = GEN_368[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_369 = {1{$random}};
  mem_reg_btb_hit = GEN_369[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_370 = {1{$random}};
  mem_reg_btb_resp_taken = GEN_370[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_371 = {1{$random}};
  mem_reg_btb_resp_mask = GEN_371[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_372 = {1{$random}};
  mem_reg_btb_resp_bridx = GEN_372[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_373 = {2{$random}};
  mem_reg_btb_resp_target = GEN_373[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_374 = {1{$random}};
  mem_reg_btb_resp_entry = GEN_374[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_375 = {1{$random}};
  mem_reg_btb_resp_bht_history = GEN_375[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_376 = {1{$random}};
  mem_reg_btb_resp_bht_value = GEN_376[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_377 = {1{$random}};
  mem_reg_xcpt = GEN_377[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_378 = {1{$random}};
  mem_reg_replay = GEN_378[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_379 = {1{$random}};
  mem_reg_flush_pipe = GEN_379[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_380 = {2{$random}};
  mem_reg_cause = GEN_380[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_381 = {1{$random}};
  mem_reg_slow_bypass = GEN_381[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_382 = {1{$random}};
  mem_reg_load = GEN_382[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_383 = {1{$random}};
  mem_reg_store = GEN_383[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_384 = {2{$random}};
  mem_reg_pc = GEN_384[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_385 = {1{$random}};
  mem_reg_inst = GEN_385[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_386 = {2{$random}};
  mem_reg_wdata = GEN_386[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_387 = {2{$random}};
  mem_reg_rs2 = GEN_387[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_388 = {1{$random}};
  wb_reg_valid = GEN_388[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_389 = {1{$random}};
  wb_reg_xcpt = GEN_389[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_390 = {1{$random}};
  wb_reg_replay = GEN_390[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_391 = {2{$random}};
  wb_reg_cause = GEN_391[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_392 = {2{$random}};
  wb_reg_pc = GEN_392[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_393 = {1{$random}};
  wb_reg_inst = GEN_393[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_394 = {2{$random}};
  wb_reg_wdata = GEN_394[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_395 = {2{$random}};
  wb_reg_rs2 = GEN_395[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_396 = {1{$random}};
  id_reg_fence = GEN_396[0:0];
  `endif
  GEN_397 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    T_7192[initvar] = GEN_397[63:0];
  `endif
  GEN_398 = {2{$random}};
  GEN_399 = {2{$random}};
  `ifdef RANDOMIZE_REG_INIT
  GEN_400 = {1{$random}};
  ex_reg_rs_bypass_0 = GEN_400[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_401 = {1{$random}};
  ex_reg_rs_bypass_1 = GEN_401[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_402 = {1{$random}};
  ex_reg_rs_lsb_0 = GEN_402[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_403 = {1{$random}};
  ex_reg_rs_lsb_1 = GEN_403[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_404 = {2{$random}};
  ex_reg_rs_msb_0 = GEN_404[61:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_405 = {2{$random}};
  ex_reg_rs_msb_1 = GEN_405[61:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_406 = {1{$random}};
  T_7896 = GEN_406[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_407 = {1{$random}};
  T_7983 = GEN_407[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_408 = {1{$random}};
  dcache_blocked = GEN_408[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_409 = {1{$random}};
  rocc_blocked = GEN_409[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_410 = {2{$random}};
  T_8257 = GEN_410[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_411 = {2{$random}};
  T_8258 = GEN_411[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_412 = {2{$random}};
  T_8260 = GEN_412[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_413 = {2{$random}};
  T_8261 = GEN_413[63:0];
  `endif
  GEN_414 = {1{$random}};
  GEN_415 = {2{$random}};
  GEN_416 = {1{$random}};
  GEN_417 = {1{$random}};
  GEN_418 = {1{$random}};
  GEN_419 = {1{$random}};
  GEN_420 = {1{$random}};
  GEN_421 = {1{$random}};
  GEN_422 = {1{$random}};
  GEN_423 = {1{$random}};
  GEN_424 = {1{$random}};
  GEN_425 = {1{$random}};
  GEN_426 = {1{$random}};
  GEN_427 = {1{$random}};
  GEN_428 = {1{$random}};
  GEN_429 = {1{$random}};
  GEN_430 = {1{$random}};
  GEN_431 = {1{$random}};
  GEN_432 = {1{$random}};
  GEN_433 = {1{$random}};
  GEN_434 = {1{$random}};
  GEN_435 = {1{$random}};
  GEN_436 = {3{$random}};
  GEN_437 = {3{$random}};
  GEN_438 = {3{$random}};
  GEN_439 = {1{$random}};
  GEN_440 = {1{$random}};
  GEN_441 = {1{$random}};
  GEN_442 = {1{$random}};
  GEN_443 = {1{$random}};
  GEN_444 = {2{$random}};
  GEN_445 = {1{$random}};
  GEN_446 = {1{$random}};
  GEN_447 = {1{$random}};
  GEN_448 = {2{$random}};
  GEN_449 = {1{$random}};
  GEN_450 = {1{$random}};
  GEN_451 = {2{$random}};
  GEN_452 = {2{$random}};
  GEN_453 = {1{$random}};
  GEN_454 = {1{$random}};
  GEN_455 = {1{$random}};
  GEN_456 = {1{$random}};
  GEN_457 = {1{$random}};
  GEN_458 = {1{$random}};
  GEN_459 = {1{$random}};
  GEN_460 = {1{$random}};
  GEN_461 = {1{$random}};
  GEN_462 = {1{$random}};
  GEN_463 = {1{$random}};
  GEN_464 = {1{$random}};
  GEN_465 = {1{$random}};
  GEN_466 = {2{$random}};
  GEN_467 = {1{$random}};
  GEN_468 = {1{$random}};
  GEN_469 = {3{$random}};
  GEN_470 = {1{$random}};
  GEN_471 = {1{$random}};
  GEN_472 = {1{$random}};
  GEN_473 = {1{$random}};
  GEN_474 = {2{$random}};
  GEN_475 = {1{$random}};
  GEN_476 = {2{$random}};
  GEN_477 = {1{$random}};
  GEN_478 = {1{$random}};
  GEN_479 = {1{$random}};
  GEN_480 = {1{$random}};
  GEN_481 = {2{$random}};
  GEN_482 = {1{$random}};
  GEN_483 = {2{$random}};
  GEN_484 = {1{$random}};
  GEN_485 = {1{$random}};
  GEN_486 = {1{$random}};
  GEN_487 = {1{$random}};
  GEN_488 = {1{$random}};
  GEN_489 = {1{$random}};
  GEN_490 = {1{$random}};
  GEN_491 = {1{$random}};
  GEN_492 = {1{$random}};
  GEN_493 = {2{$random}};
  GEN_494 = {1{$random}};
  GEN_495 = {1{$random}};
  GEN_496 = {1{$random}};
  GEN_497 = {1{$random}};
  GEN_498 = {1{$random}};
  GEN_499 = {1{$random}};
  GEN_500 = {1{$random}};
  GEN_501 = {1{$random}};
  GEN_502 = {1{$random}};
  GEN_503 = {1{$random}};
  GEN_504 = {1{$random}};
  GEN_505 = {1{$random}};
  GEN_506 = {1{$random}};
  GEN_507 = {1{$random}};
  GEN_508 = {1{$random}};
  GEN_509 = {1{$random}};
  GEN_510 = {1{$random}};
  GEN_511 = {1{$random}};
  GEN_512 = {1{$random}};
  GEN_513 = {1{$random}};
  GEN_514 = {1{$random}};
  GEN_515 = {3{$random}};
  GEN_516 = {3{$random}};
  GEN_517 = {3{$random}};
  GEN_518 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_legal <= id_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_fp <= id_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_rocc <= id_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_branch <= id_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_jal <= id_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_jalr <= id_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_rxs2 <= id_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_rxs1 <= id_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(id_xcpt) begin
          if(T_7562) begin
            ex_ctrl_sel_alu2 <= 2'h1;
          end else begin
            ex_ctrl_sel_alu2 <= 2'h0;
          end
        end else begin
          ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(id_xcpt) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else begin
          ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_sel_imm <= id_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(id_xcpt) begin
          ex_ctrl_alu_dw <= 1'h1;
        end else begin
          ex_ctrl_alu_dw <= id_ctrl_alu_dw;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(id_xcpt) begin
          ex_ctrl_alu_fn <= 4'h0;
        end else begin
          ex_ctrl_alu_fn <= id_ctrl_alu_fn;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_mem <= id_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_mem_type <= id_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_rfs1 <= id_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_rfs2 <= id_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_rfs3 <= id_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_wfd <= id_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_div <= id_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_wxd <= id_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(id_csr_ren) begin
          ex_ctrl_csr <= 3'h5;
        end else begin
          ex_ctrl_csr <= id_ctrl_csr;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(T_7566) begin
          ex_ctrl_fence_i <= 1'h1;
        end else begin
          ex_ctrl_fence_i <= id_ctrl_fence_i;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_fence <= id_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_ctrl_amo <= id_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_legal <= ex_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fp <= ex_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rocc <= ex_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_branch <= ex_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_jal <= ex_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_jalr <= ex_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rxs2 <= ex_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rxs1 <= ex_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_alu2 <= ex_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_alu1 <= ex_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_imm <= ex_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_alu_dw <= ex_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_alu_fn <= ex_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem <= ex_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem_cmd <= ex_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem_type <= ex_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs1 <= ex_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs2 <= ex_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs3 <= ex_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_wfd <= ex_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_div <= ex_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_wxd <= ex_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_csr <= ex_ctrl_csr;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fence_i <= ex_ctrl_fence_i;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fence <= ex_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_amo <= ex_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_legal <= mem_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_fp <= mem_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_rocc <= mem_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_branch <= mem_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_jal <= mem_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_jalr <= mem_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_rxs2 <= mem_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_rxs1 <= mem_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_sel_alu2 <= mem_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_sel_alu1 <= mem_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_sel_imm <= mem_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_alu_dw <= mem_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_alu_fn <= mem_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_mem <= mem_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_mem_cmd <= mem_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_mem_type <= mem_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_rfs1 <= mem_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_rfs2 <= mem_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_rfs3 <= mem_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_wfd <= mem_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_div <= mem_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_wxd <= mem_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_csr <= mem_ctrl_csr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_fence_i <= mem_ctrl_fence_i;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_fence <= mem_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_ctrl_amo <= mem_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt_interrupt <= T_7554;
    end
    if(1'h0) begin
    end else begin
      ex_reg_valid <= T_7543;
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(id_xcpt) begin
          if(T_7562) begin
            ex_reg_rvc <= 1'h1;
          end else begin
            ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
          end
        end else begin
          ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
        end
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_hit <= ibuf_io_inst_0_bits_btb_hit;
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_taken <= ibuf_io_btb_resp_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_mask <= ibuf_io_btb_resp_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_bridx <= ibuf_io_btb_resp_bridx;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_target <= ibuf_io_btb_resp_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_entry <= ibuf_io_btb_resp_entry;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_bht_history <= ibuf_io_btb_resp_bht_history;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_bht_value <= ibuf_io_btb_resp_bht_value;
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt <= T_7550;
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(T_7566) begin
          ex_reg_flush_pipe <= 1'h1;
        end else begin
          ex_reg_flush_pipe <= T_7565;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_reg_load_use <= id_load_use;
      end
    end
    if(1'h0) begin
    end else begin
      if(id_xcpt) begin
        if(csr_io_interrupt) begin
          ex_reg_cause <= csr_io_interrupt_cause;
        end else begin
          ex_reg_cause <= {{60'd0}, T_7407};
        end
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_replay <= T_7547;
    end
    if(1'h0) begin
    end else begin
      if(T_7602) begin
        ex_reg_pc <= ibuf_io_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7602) begin
        ex_reg_inst <= ibuf_io_inst_0_bits_inst_bits;
      end
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt_interrupt <= T_7840;
    end
    if(1'h0) begin
    end else begin
      mem_reg_valid <= T_7831;
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_rvc <= ex_reg_rvc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_btb_hit <= ex_reg_btb_hit;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_mask <= ex_reg_btb_resp_mask;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bridx <= ex_reg_btb_resp_bridx;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
        end
      end
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt <= T_7837;
    end
    if(1'h0) begin
    end else begin
      mem_reg_replay <= T_7834;
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_flush_pipe <= ex_reg_flush_pipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_xcpt) begin
        if(T_7634) begin
          mem_reg_cause <= ex_reg_cause;
        end else begin
          mem_reg_cause <= 64'h2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_slow_bypass <= ex_slow_bypass;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_load <= T_7850;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_store <= T_7858;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_pc <= ex_reg_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_inst <= ex_reg_inst;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_wdata <= alu_io_out;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(T_7860) begin
          if(ex_reg_rs_bypass_1) begin
            mem_reg_rs2 <= GEN_1;
          end else begin
            mem_reg_rs2 <= T_7453;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      wb_reg_valid <= T_7900;
    end
    if(1'h0) begin
    end else begin
      wb_reg_xcpt <= T_7906;
    end
    if(1'h0) begin
    end else begin
      wb_reg_replay <= T_7903;
    end
    if(1'h0) begin
    end else begin
      if(mem_xcpt) begin
        if(T_7886) begin
          wb_reg_cause <= mem_reg_cause;
        end else begin
          wb_reg_cause <= {{60'd0}, mem_new_cause};
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_reg_pc <= mem_reg_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        wb_reg_inst <= mem_reg_inst;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        if(T_7912) begin
          wb_reg_wdata <= io_fpu_toint_data;
        end else begin
          wb_reg_wdata <= mem_int_wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7908) begin
        if(mem_ctrl_rocc) begin
          wb_reg_rs2 <= mem_reg_rs2;
        end
      end
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T_7389;
    end
    if(T_7192_T_7944_en & T_7192_T_7944_mask) begin
      T_7192[T_7192_T_7944_addr] <= T_7192_T_7944_data;
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_reg_rs_bypass_0 <= T_7571;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        ex_reg_rs_bypass_1 <= T_7586;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(T_7581) begin
          ex_reg_rs_lsb_0 <= T_7582;
        end else begin
          if(T_7417) begin
            ex_reg_rs_lsb_0 <= 2'h0;
          end else begin
            if(id_bypass_src_0_1) begin
              ex_reg_rs_lsb_0 <= 2'h1;
            end else begin
              if(id_bypass_src_0_2) begin
                ex_reg_rs_lsb_0 <= 2'h2;
              end else begin
                ex_reg_rs_lsb_0 <= 2'h3;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(T_7596) begin
          ex_reg_rs_lsb_1 <= T_7597;
        end else begin
          if(T_7421) begin
            ex_reg_rs_lsb_1 <= 2'h0;
          end else begin
            if(id_bypass_src_1_1) begin
              ex_reg_rs_lsb_1 <= 2'h1;
            end else begin
              if(id_bypass_src_1_2) begin
                ex_reg_rs_lsb_1 <= 2'h2;
              end else begin
                ex_reg_rs_lsb_1 <= 2'h3;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(T_7581) begin
          ex_reg_rs_msb_0 <= T_7583;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7543) begin
        if(T_7596) begin
          ex_reg_rs_msb_1 <= T_7598;
        end
      end
    end
    if(1'h0) begin
    end else begin
      T_7896 <= T_7895;
    end
    if(reset) begin
      T_7983 <= 32'h0;
    end else begin
      if(T_8010) begin
        T_7983 <= T_8009;
      end else begin
        if(ll_wen) begin
          T_7983 <= T_7992;
        end
      end
    end
    if(1'h0) begin
    end else begin
      dcache_blocked <= T_8091;
    end
    if(1'h0) begin
    end else begin
      rocc_blocked <= T_8099;
    end
    if(1'h0) begin
    end else begin
      if(ex_reg_rs_bypass_0) begin
        T_8257 <= GEN_0;
      end else begin
        T_8257 <= T_7452;
      end
    end
    if(1'h0) begin
    end else begin
      T_8258 <= T_8257;
    end
    if(1'h0) begin
    end else begin
      if(ex_reg_rs_bypass_1) begin
        T_8260 <= GEN_1;
      end else begin
        T_8260 <= T_7453;
      end
    end
    if(1'h0) begin
    end else begin
      T_8261 <= T_8260;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_8200 & T_8208) begin
          $fwrite(32'h80000002,"Assertion failed\n    at rocket.scala:632 assert(io.dmem.xcpt.asUInt.orR) // make sure s1_kill is exhaustive\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_8200 & T_8208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_8263) begin
          $fwrite(32'h80000002,"C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n",io_prci_id,T_8253,wb_valid,wb_reg_pc,T_8255,rf_wdata,rf_wen,T_8256,T_8258,T_8259,T_8261,wb_reg_inst,wb_reg_inst);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module FlowThroughSerializer(
  input   clk,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input  [2:0] io_in_bits_addr_beat,
  input   io_in_bits_client_xact_id,
  input  [1:0] io_in_bits_manager_xact_id,
  input   io_in_bits_is_builtin_type,
  input  [3:0] io_in_bits_g_type,
  input  [63:0] io_in_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_client_xact_id,
  output [1:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_cnt,
  output  io_done
);
  assign io_in_ready = io_out_ready;
  assign io_out_valid = io_in_valid;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_data = io_in_bits_data;
  assign io_cnt = 1'h0;
  assign io_done = 1'h1;
endmodule
module ICache(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [38:0] io_req_bits_addr,
  input  [19:0] io_s1_ppn,
  input   io_s1_kill,
  input   io_s2_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [15:0] io_resp_bits_data,
  output [63:0] io_resp_bits_datablock,
  input   io_invalidate,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output  io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [10:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input   io_mem_grant_bits_client_xact_id,
  input  [1:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
  reg [1:0] state;
  reg [31:0] GEN_4;
  reg  invalidated;
  reg [31:0] GEN_5;
  wire  stall;
  wire  rdy;
  reg [31:0] refill_addr;
  reg [31:0] GEN_6;
  wire  s1_any_tag_hit;
  reg  s1_valid;
  reg [31:0] GEN_7;
  reg [38:0] s1_vaddr;
  reg [63:0] GEN_8;
  wire [11:0] T_827;
  wire [31:0] s1_paddr;
  wire [19:0] s1_tag;
  wire  T_828;
  wire  s0_valid;
  wire [38:0] s0_vaddr;
  wire  T_830;
  wire  T_833;
  wire  T_834;
  wire  T_835;
  wire [38:0] GEN_0;
  wire  T_839;
  wire  T_840;
  wire  out_valid;
  wire [5:0] s1_idx;
  wire  s1_hit;
  wire  T_842;
  wire  s1_miss;
  wire  T_845;
  wire  T_846;
  wire  T_848;
  wire [31:0] GEN_1;
  wire [19:0] refill_tag;
  wire  FlowThroughSerializer_1_clk;
  wire  FlowThroughSerializer_1_reset;
  wire  FlowThroughSerializer_1_io_in_ready;
  wire  FlowThroughSerializer_1_io_in_valid;
  wire [2:0] FlowThroughSerializer_1_io_in_bits_addr_beat;
  wire  FlowThroughSerializer_1_io_in_bits_client_xact_id;
  wire [1:0] FlowThroughSerializer_1_io_in_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_io_in_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_io_in_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_io_in_bits_data;
  wire  FlowThroughSerializer_1_io_out_ready;
  wire  FlowThroughSerializer_1_io_out_valid;
  wire [2:0] FlowThroughSerializer_1_io_out_bits_addr_beat;
  wire  FlowThroughSerializer_1_io_out_bits_client_xact_id;
  wire [1:0] FlowThroughSerializer_1_io_out_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_io_out_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_io_out_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_io_out_bits_data;
  wire  FlowThroughSerializer_1_io_cnt;
  wire  FlowThroughSerializer_1_io_done;
  wire  T_849;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_9;
  wire  T_852;
  wire [3:0] T_854;
  wire [2:0] T_855;
  wire [2:0] GEN_2;
  wire  refill_wrap;
  wire  T_856;
  wire  refill_done;
  reg [19:0] tag_array_0 [0:63];
  reg [31:0] GEN_10;
  wire [19:0] tag_array_0_tag_rdata_data;
  wire [5:0] tag_array_0_tag_rdata_addr;
  wire  tag_array_0_tag_rdata_en;
  reg [5:0] GEN_11;
  reg [31:0] GEN_12;
  wire [19:0] tag_array_0_T_893_data;
  wire [5:0] tag_array_0_T_893_addr;
  wire  tag_array_0_T_893_mask;
  wire  tag_array_0_T_893_en;
  wire [5:0] T_866;
  wire  T_868;
  wire  T_869;
  wire [5:0] T_871;
  wire [19:0] T_880_0;
  wire  T_889_0;
  wire  GEN_13;
  reg [63:0] vb_array;
  reg [63:0] GEN_18;
  wire  T_897;
  wire  T_898;
  wire [6:0] T_899;
  wire [127:0] T_902;
  wire [127:0] GEN_38;
  wire [127:0] T_903;
  wire [63:0] T_904;
  wire [127:0] GEN_39;
  wire [127:0] T_905;
  wire [127:0] T_906;
  wire [127:0] GEN_14;
  wire [127:0] GEN_15;
  wire  GEN_16;
  wire  s1_disparity_0;
  wire  T_917;
  wire [127:0] GEN_17;
  wire  s1_tag_match_0;
  wire  s1_tag_hit_0;
  wire [63:0] s1_dout_0;
  wire  T_950;
  wire [63:0] T_954;
  wire  T_955;
  wire  T_957;
  wire [19:0] T_961;
  wire  T_962;
  wire  T_963;
  wire  T_970;
  wire  T_971;
  reg [63:0] T_974 [0:511];
  reg [63:0] GEN_19;
  wire [63:0] T_974_T_987_data;
  wire [8:0] T_974_T_987_addr;
  wire  T_974_T_987_en;
  reg [8:0] GEN_20;
  reg [31:0] GEN_22;
  wire [63:0] T_974_T_980_data;
  wire [8:0] T_974_T_980_addr;
  wire  T_974_T_980_mask;
  wire  T_974_T_980_en;
  wire  T_977;
  wire [8:0] GEN_42;
  wire [8:0] T_978;
  wire [8:0] GEN_43;
  wire [8:0] T_979;
  wire [63:0] GEN_21;
  wire [8:0] T_981;
  wire  T_983;
  wire  T_984;
  wire [8:0] T_986;
  wire  T_989;
  reg  T_990;
  reg [31:0] GEN_23;
  wire  GEN_25;
  reg  T_995_0;
  reg [31:0] GEN_24;
  wire  GEN_26;
  reg [63:0] T_1001_0;
  reg [63:0] GEN_40;
  wire [63:0] GEN_27;
  wire  T_1003;
  wire  T_1005;
  wire  T_1006;
  wire [25:0] T_1007;
  wire [25:0] T_1131_addr_block;
  wire  T_1131_client_xact_id;
  wire [2:0] T_1131_addr_beat;
  wire  T_1131_is_builtin_type;
  wire [2:0] T_1131_a_type;
  wire [10:0] T_1131_union;
  wire [63:0] T_1131_data;
  wire  T_1159;
  wire [1:0] GEN_28;
  wire [1:0] GEN_29;
  wire  GEN_30;
  wire  T_1161;
  wire [1:0] GEN_31;
  wire [1:0] GEN_32;
  wire [1:0] GEN_33;
  wire  T_1162;
  wire [1:0] GEN_34;
  wire [1:0] GEN_35;
  wire  T_1163;
  wire [1:0] GEN_36;
  wire [1:0] GEN_37;
  wire [15:0] GEN_3;
  reg [31:0] GEN_41;
  FlowThroughSerializer FlowThroughSerializer_1 (
    .clk(FlowThroughSerializer_1_clk),
    .reset(FlowThroughSerializer_1_reset),
    .io_in_ready(FlowThroughSerializer_1_io_in_ready),
    .io_in_valid(FlowThroughSerializer_1_io_in_valid),
    .io_in_bits_addr_beat(FlowThroughSerializer_1_io_in_bits_addr_beat),
    .io_in_bits_client_xact_id(FlowThroughSerializer_1_io_in_bits_client_xact_id),
    .io_in_bits_manager_xact_id(FlowThroughSerializer_1_io_in_bits_manager_xact_id),
    .io_in_bits_is_builtin_type(FlowThroughSerializer_1_io_in_bits_is_builtin_type),
    .io_in_bits_g_type(FlowThroughSerializer_1_io_in_bits_g_type),
    .io_in_bits_data(FlowThroughSerializer_1_io_in_bits_data),
    .io_out_ready(FlowThroughSerializer_1_io_out_ready),
    .io_out_valid(FlowThroughSerializer_1_io_out_valid),
    .io_out_bits_addr_beat(FlowThroughSerializer_1_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(FlowThroughSerializer_1_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(FlowThroughSerializer_1_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(FlowThroughSerializer_1_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(FlowThroughSerializer_1_io_out_bits_g_type),
    .io_out_bits_data(FlowThroughSerializer_1_io_out_bits_data),
    .io_cnt(FlowThroughSerializer_1_io_cnt),
    .io_done(FlowThroughSerializer_1_io_done)
  );
  assign io_resp_valid = T_990;
  assign io_resp_bits_data = GEN_3;
  assign io_resp_bits_datablock = T_1001_0;
  assign io_mem_acquire_valid = T_1006;
  assign io_mem_acquire_bits_addr_block = T_1131_addr_block;
  assign io_mem_acquire_bits_client_xact_id = T_1131_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = T_1131_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = T_1131_is_builtin_type;
  assign io_mem_acquire_bits_a_type = T_1131_a_type;
  assign io_mem_acquire_bits_union = T_1131_union;
  assign io_mem_acquire_bits_data = T_1131_data;
  assign io_mem_grant_ready = FlowThroughSerializer_1_io_in_ready;
  assign stall = io_resp_ready == 1'h0;
  assign rdy = T_846;
  assign s1_any_tag_hit = T_971;
  assign T_827 = s1_vaddr[11:0];
  assign s1_paddr = {io_s1_ppn,T_827};
  assign s1_tag = s1_paddr[31:12];
  assign T_828 = s1_valid & stall;
  assign s0_valid = io_req_valid | T_828;
  assign s0_vaddr = T_828 ? s1_vaddr : io_req_bits_addr;
  assign T_830 = io_req_valid & rdy;
  assign T_833 = io_s1_kill == 1'h0;
  assign T_834 = T_828 & T_833;
  assign T_835 = T_830 | T_834;
  assign GEN_0 = T_830 ? io_req_bits_addr : s1_vaddr;
  assign T_839 = s1_valid & T_833;
  assign T_840 = state == 2'h0;
  assign out_valid = T_839 & T_840;
  assign s1_idx = s1_vaddr[11:6];
  assign s1_hit = out_valid & s1_any_tag_hit;
  assign T_842 = s1_any_tag_hit == 1'h0;
  assign s1_miss = out_valid & T_842;
  assign T_845 = s1_miss == 1'h0;
  assign T_846 = T_840 & T_845;
  assign T_848 = s1_miss & T_840;
  assign GEN_1 = T_848 ? s1_paddr : refill_addr;
  assign refill_tag = refill_addr[31:12];
  assign FlowThroughSerializer_1_clk = clk;
  assign FlowThroughSerializer_1_reset = reset;
  assign FlowThroughSerializer_1_io_in_valid = io_mem_grant_valid;
  assign FlowThroughSerializer_1_io_in_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign FlowThroughSerializer_1_io_in_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign FlowThroughSerializer_1_io_in_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign FlowThroughSerializer_1_io_in_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign FlowThroughSerializer_1_io_in_bits_g_type = io_mem_grant_bits_g_type;
  assign FlowThroughSerializer_1_io_in_bits_data = io_mem_grant_bits_data;
  assign FlowThroughSerializer_1_io_out_ready = 1'h1;
  assign T_849 = FlowThroughSerializer_1_io_out_ready & FlowThroughSerializer_1_io_out_valid;
  assign T_852 = refill_cnt == 3'h7;
  assign T_854 = refill_cnt + 3'h1;
  assign T_855 = T_854[2:0];
  assign GEN_2 = T_849 ? T_855 : refill_cnt;
  assign refill_wrap = T_849 & T_852;
  assign T_856 = state == 2'h3;
  assign refill_done = T_856 & refill_wrap;
  assign tag_array_0_tag_rdata_addr = T_871;
  assign tag_array_0_tag_rdata_en = T_869;
  assign tag_array_0_tag_rdata_data = tag_array_0[GEN_11];
  assign tag_array_0_T_893_data = T_880_0;
  assign tag_array_0_T_893_addr = s1_idx;
  assign tag_array_0_T_893_mask = GEN_13;
  assign tag_array_0_T_893_en = refill_done;
  assign T_866 = s0_vaddr[11:6];
  assign T_868 = refill_done == 1'h0;
  assign T_869 = T_868 & s0_valid;
  assign T_871 = T_866;
  assign T_880_0 = refill_tag;
  assign T_889_0 = 1'h1;
  assign GEN_13 = refill_done ? T_889_0 : 1'h0;
  assign T_897 = invalidated == 1'h0;
  assign T_898 = refill_done & T_897;
  assign T_899 = {1'h0,s1_idx};
  assign T_902 = 128'h1 << T_899;
  assign GEN_38 = {{64'd0}, vb_array};
  assign T_903 = GEN_38 | T_902;
  assign T_904 = ~ vb_array;
  assign GEN_39 = {{64'd0}, T_904};
  assign T_905 = GEN_39 | T_902;
  assign T_906 = ~ T_905;
  assign GEN_14 = T_898 ? T_903 : {{64'd0}, vb_array};
  assign GEN_15 = io_invalidate ? 128'h0 : GEN_14;
  assign GEN_16 = io_invalidate ? 1'h1 : invalidated;
  assign s1_disparity_0 = 1'h0;
  assign T_917 = s1_valid & s1_disparity_0;
  assign GEN_17 = T_917 ? T_906 : GEN_15;
  assign s1_tag_match_0 = T_962;
  assign s1_tag_hit_0 = T_963;
  assign s1_dout_0 = T_974_T_987_data;
  assign T_950 = io_invalidate == 1'h0;
  assign T_954 = vb_array >> T_899;
  assign T_955 = T_954[0];
  assign T_957 = T_950 & T_955;
  assign T_961 = tag_array_0_tag_rdata_data;
  assign T_962 = T_961 == s1_tag;
  assign T_963 = T_957 & s1_tag_match_0;
  assign T_970 = s1_disparity_0 == 1'h0;
  assign T_971 = s1_tag_hit_0 & T_970;
  assign T_974_T_987_addr = T_986;
  assign T_974_T_987_en = T_984;
  assign T_974_T_987_data = T_974[GEN_20];
  assign T_974_T_980_data = GEN_21;
  assign T_974_T_980_addr = T_979;
  assign T_974_T_980_mask = T_977;
  assign T_974_T_980_en = T_977;
  assign T_977 = FlowThroughSerializer_1_io_out_valid;
  assign GEN_42 = {{3'd0}, s1_idx};
  assign T_978 = GEN_42 << 3;
  assign GEN_43 = {{6'd0}, refill_cnt};
  assign T_979 = T_978 | GEN_43;
  assign GEN_21 = FlowThroughSerializer_1_io_out_bits_data;
  assign T_981 = s0_vaddr[11:3];
  assign T_983 = T_977 == 1'h0;
  assign T_984 = T_983 & s0_valid;
  assign T_986 = T_981;
  assign T_989 = stall == 1'h0;
  assign GEN_25 = T_989 ? s1_hit : T_990;
  assign GEN_26 = T_989 ? s1_tag_hit_0 : T_995_0;
  assign GEN_27 = T_989 ? s1_dout_0 : T_1001_0;
  assign T_1003 = state == 2'h1;
  assign T_1005 = io_s2_kill == 1'h0;
  assign T_1006 = T_1003 & T_1005;
  assign T_1007 = refill_addr[31:6];
  assign T_1131_addr_block = T_1007;
  assign T_1131_client_xact_id = 1'h0;
  assign T_1131_addr_beat = 3'h0;
  assign T_1131_is_builtin_type = 1'h1;
  assign T_1131_a_type = 3'h1;
  assign T_1131_union = 11'hc1;
  assign T_1131_data = 64'h0;
  assign T_1159 = 2'h0 == state;
  assign GEN_28 = s1_miss ? 2'h1 : state;
  assign GEN_29 = T_1159 ? GEN_28 : state;
  assign GEN_30 = T_1159 ? 1'h0 : GEN_16;
  assign T_1161 = 2'h1 == state;
  assign GEN_31 = io_mem_acquire_ready ? 2'h2 : GEN_29;
  assign GEN_32 = io_s2_kill ? 2'h0 : GEN_31;
  assign GEN_33 = T_1161 ? GEN_32 : GEN_29;
  assign T_1162 = 2'h2 == state;
  assign GEN_34 = io_mem_grant_valid ? 2'h3 : GEN_33;
  assign GEN_35 = T_1162 ? GEN_34 : GEN_33;
  assign T_1163 = 2'h3 == state;
  assign GEN_36 = refill_done ? 2'h0 : GEN_35;
  assign GEN_37 = T_1163 ? GEN_36 : GEN_35;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_41[15:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {1{$random}};
  state = GEN_4[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  invalidated = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  refill_addr = GEN_6[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  s1_valid = GEN_7[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {2{$random}};
  s1_vaddr = GEN_8[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {1{$random}};
  refill_cnt = GEN_9[2:0];
  `endif
  GEN_10 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = GEN_10[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_12 = {1{$random}};
  GEN_11 = GEN_12[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {2{$random}};
  vb_array = GEN_18[63:0];
  `endif
  GEN_19 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_974[initvar] = GEN_19[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_22 = {1{$random}};
  GEN_20 = GEN_22[8:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_23 = {1{$random}};
  T_990 = GEN_23[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_24 = {1{$random}};
  T_995_0 = GEN_24[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {2{$random}};
  T_1001_0 = GEN_40[63:0];
  `endif
  GEN_41 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else begin
      if(T_1163) begin
        if(refill_done) begin
          state <= 2'h0;
        end else begin
          if(T_1162) begin
            if(io_mem_grant_valid) begin
              state <= 2'h3;
            end else begin
              if(T_1161) begin
                if(io_s2_kill) begin
                  state <= 2'h0;
                end else begin
                  if(io_mem_acquire_ready) begin
                    state <= 2'h2;
                  end else begin
                    if(T_1159) begin
                      if(s1_miss) begin
                        state <= 2'h1;
                      end
                    end
                  end
                end
              end else begin
                if(T_1159) begin
                  if(s1_miss) begin
                    state <= 2'h1;
                  end
                end
              end
            end
          end else begin
            if(T_1161) begin
              if(io_s2_kill) begin
                state <= 2'h0;
              end else begin
                if(io_mem_acquire_ready) begin
                  state <= 2'h2;
                end else begin
                  if(T_1159) begin
                    if(s1_miss) begin
                      state <= 2'h1;
                    end
                  end
                end
              end
            end else begin
              if(T_1159) begin
                if(s1_miss) begin
                  state <= 2'h1;
                end
              end
            end
          end
        end
      end else begin
        if(T_1162) begin
          if(io_mem_grant_valid) begin
            state <= 2'h3;
          end else begin
            if(T_1161) begin
              if(io_s2_kill) begin
                state <= 2'h0;
              end else begin
                if(io_mem_acquire_ready) begin
                  state <= 2'h2;
                end else begin
                  state <= GEN_29;
                end
              end
            end else begin
              state <= GEN_29;
            end
          end
        end else begin
          if(T_1161) begin
            if(io_s2_kill) begin
              state <= 2'h0;
            end else begin
              if(io_mem_acquire_ready) begin
                state <= 2'h2;
              end else begin
                state <= GEN_29;
              end
            end
          end else begin
            state <= GEN_29;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1159) begin
        invalidated <= 1'h0;
      end else begin
        if(io_invalidate) begin
          invalidated <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_848) begin
        refill_addr <= s1_paddr;
      end
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_835;
    end
    if(1'h0) begin
    end else begin
      if(T_830) begin
        s1_vaddr <= io_req_bits_addr;
      end
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      if(T_849) begin
        refill_cnt <= T_855;
      end
    end
    if(tag_array_0_tag_rdata_en) begin
      GEN_11 <= tag_array_0_tag_rdata_addr;
    end
    if(tag_array_0_T_893_en & tag_array_0_T_893_mask) begin
      tag_array_0[tag_array_0_T_893_addr] <= tag_array_0_T_893_data;
    end
    if(reset) begin
      vb_array <= 64'h0;
    end else begin
      vb_array <= GEN_17[63:0];
    end
    if(T_974_T_987_en) begin
      GEN_20 <= T_974_T_987_addr;
    end
    if(T_974_T_980_en & T_974_T_980_mask) begin
      T_974[T_974_T_980_addr] <= T_974_T_980_data;
    end
    if(1'h0) begin
    end else begin
      if(T_989) begin
        T_990 <= s1_hit;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_989) begin
        T_995_0 <= s1_tag_hit_0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_989) begin
        T_1001_0 <= s1_dout_0;
      end
    end
  end
endmodule
module TLB(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [27:0] io_req_bits_vpn,
  input   io_req_bits_passthrough,
  input   io_req_bits_instruction,
  input   io_req_bits_store,
  output  io_resp_miss,
  output [19:0] io_resp_ppn,
  output  io_resp_xcpt_ld,
  output  io_resp_xcpt_st,
  output  io_resp_xcpt_if,
  output  io_resp_cacheable,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_pum,
  output  io_ptw_req_bits_mxr,
  output [26:0] io_ptw_req_bits_addr,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [15:0] io_ptw_resp_bits_pte_reserved_for_hardware,
  input  [37:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_a,
  input   io_ptw_resp_bits_pte_g,
  input   io_ptw_resp_bits_pte_u,
  input   io_ptw_resp_bits_pte_x,
  input   io_ptw_resp_bits_pte_w,
  input   io_ptw_resp_bits_pte_r,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [37:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [3:0] io_ptw_status_zero1,
  input   io_ptw_status_mxr,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie
);
  reg [3:0] valid;
  reg [31:0] GEN_2;
  reg [19:0] ppns_0;
  reg [31:0] GEN_3;
  reg [19:0] ppns_1;
  reg [31:0] GEN_4;
  reg [19:0] ppns_2;
  reg [31:0] GEN_5;
  reg [19:0] ppns_3;
  reg [31:0] GEN_6;
  reg [33:0] tags_0;
  reg [63:0] GEN_7;
  reg [33:0] tags_1;
  reg [63:0] GEN_8;
  reg [33:0] tags_2;
  reg [63:0] GEN_9;
  reg [33:0] tags_3;
  reg [63:0] GEN_10;
  reg [1:0] state;
  reg [31:0] GEN_11;
  reg [33:0] r_refill_tag;
  reg [63:0] GEN_12;
  reg [1:0] r_refill_waddr;
  reg [31:0] GEN_13;
  reg [27:0] r_req_vpn;
  reg [31:0] GEN_14;
  reg  r_req_passthrough;
  reg [31:0] GEN_15;
  reg  r_req_instruction;
  reg [31:0] GEN_16;
  reg  r_req_store;
  reg [31:0] GEN_17;
  wire  T_217;
  wire  do_mprv;
  wire [1:0] priv;
  wire  priv_s;
  wire [19:0] passthrough_ppn;
  wire [31:0] GEN_29;
  wire [31:0] T_224;
  wire  T_228;
  wire [2:0] T_232;
  wire  T_234;
  wire  T_236;
  wire  T_237;
  wire [2:0] T_240;
  wire  T_242;
  wire  T_244;
  wire  T_245;
  wire [2:0] T_248;
  wire  T_250;
  wire  T_252;
  wire  T_253;
  wire [2:0] T_256;
  wire  T_258;
  wire  T_260;
  wire  T_261;
  wire [2:0] T_264;
  wire [2:0] T_269;
  wire [2:0] T_270;
  wire [2:0] T_271;
  wire [2:0] T_272;
  wire  prot_x;
  wire  prot_w;
  wire  prot_r;
  wire  T_280;
  wire  T_281;
  wire  T_282;
  reg [15:0] pte_array_reserved_for_hardware;
  reg [31:0] GEN_18;
  reg [37:0] pte_array_ppn;
  reg [63:0] GEN_19;
  reg [1:0] pte_array_reserved_for_software;
  reg [31:0] GEN_20;
  reg  pte_array_d;
  reg [31:0] GEN_21;
  reg  pte_array_a;
  reg [31:0] GEN_22;
  reg  pte_array_g;
  reg [31:0] GEN_23;
  reg  pte_array_u;
  reg [31:0] GEN_24;
  reg  pte_array_x;
  reg [31:0] GEN_25;
  reg  pte_array_w;
  reg [31:0] GEN_26;
  reg  pte_array_r;
  reg [31:0] GEN_27;
  reg  pte_array_v;
  reg [31:0] GEN_30;
  reg [3:0] u_array;
  reg [31:0] GEN_31;
  reg [3:0] sw_array;
  reg [31:0] GEN_33;
  reg [3:0] sx_array;
  reg [31:0] GEN_34;
  reg [3:0] sr_array;
  reg [31:0] GEN_35;
  reg [3:0] xr_array;
  reg [31:0] GEN_36;
  reg [3:0] cash_array;
  reg [31:0] GEN_37;
  reg [3:0] dirty_array;
  reg [31:0] GEN_38;
  wire [19:0] GEN_0;
  wire [33:0] GEN_1;
  reg [3:0] T_403;
  reg [31:0] GEN_39;
  wire [3:0] T_430;
  wire [3:0] T_431;
  wire [3:0] priv_ok;
  wire [3:0] T_432;
  wire [4:0] w_array;
  wire [3:0] T_433;
  wire [4:0] x_array;
  wire [3:0] T_435;
  wire [3:0] T_436;
  wire [3:0] T_437;
  wire [4:0] r_array;
  wire [4:0] c_array;
  wire  T_438;
  wire  T_439;
  wire  bad_va;
  wire [1:0] T_467;
  wire [3:0] GEN_32;
  wire [3:0] T_468;
  wire [3:0] T_478;
  wire [3:0] T_479;
  wire [3:0] GEN_28;
  wire  T_485;
  wire [4:0] T_486;
  wire [4:0] T_487;
  wire  T_489;
  wire  T_490;
  wire [4:0] T_491;
  wire [4:0] T_492;
  wire  T_494;
  wire  T_495;
  wire [4:0] T_496;
  wire [4:0] T_497;
  wire  T_499;
  wire  T_500;
  wire [4:0] T_501;
  wire  T_503;
  wire [19:0] T_520;
  wire  T_521;
  assign io_req_ready = T_485;
  assign io_resp_miss = 1'h0;
  assign io_resp_ppn = T_520;
  assign io_resp_xcpt_ld = T_490;
  assign io_resp_xcpt_st = T_495;
  assign io_resp_xcpt_if = T_500;
  assign io_resp_cacheable = T_503;
  assign io_ptw_req_valid = T_521;
  assign io_ptw_req_bits_prv = io_ptw_status_prv;
  assign io_ptw_req_bits_pum = io_ptw_status_pum;
  assign io_ptw_req_bits_mxr = io_ptw_status_mxr;
  assign io_ptw_req_bits_addr = r_refill_tag[26:0];
  assign io_ptw_req_bits_store = r_req_store;
  assign io_ptw_req_bits_fetch = r_req_instruction;
  assign T_217 = io_req_bits_instruction == 1'h0;
  assign do_mprv = io_ptw_status_mprv & T_217;
  assign priv = do_mprv ? io_ptw_status_mpp : io_ptw_status_prv;
  assign priv_s = priv == 2'h1;
  assign passthrough_ppn = io_req_bits_vpn[19:0];
  assign GEN_29 = {{12'd0}, passthrough_ppn};
  assign T_224 = GEN_29 << 12;
  assign T_228 = T_224 < 32'h1000;
  assign T_232 = T_228 ? 3'h7 : 3'h0;
  assign T_234 = 32'h1000 <= T_224;
  assign T_236 = T_224 < 32'h2000;
  assign T_237 = T_234 & T_236;
  assign T_240 = T_237 ? 3'h5 : 3'h0;
  assign T_242 = 32'h40000000 <= T_224;
  assign T_244 = T_224 < 32'h44000000;
  assign T_245 = T_242 & T_244;
  assign T_248 = T_245 ? 3'h3 : 3'h0;
  assign T_250 = 32'h44000000 <= T_224;
  assign T_252 = T_224 < 32'h48000000;
  assign T_253 = T_250 & T_252;
  assign T_256 = T_253 ? 3'h3 : 3'h0;
  assign T_258 = 32'h80000000 <= T_224;
  assign T_260 = T_224 < 32'h90000000;
  assign T_261 = T_258 & T_260;
  assign T_264 = T_261 ? 3'h7 : 3'h0;
  assign T_269 = T_232 | T_240;
  assign T_270 = T_269 | T_248;
  assign T_271 = T_270 | T_256;
  assign T_272 = T_271 | T_264;
  assign prot_x = T_282;
  assign prot_w = T_281;
  assign prot_r = T_280;
  assign T_280 = T_272[0];
  assign T_281 = T_272[1];
  assign T_282 = T_272[2];
  assign GEN_0 = io_ptw_resp_bits_pte_ppn[19:0];
  assign GEN_1 = r_refill_tag;
  assign T_430 = io_ptw_status_pum ? u_array : 4'h0;
  assign T_431 = ~ T_430;
  assign priv_ok = priv_s ? T_431 : u_array;
  assign T_432 = priv_ok & sw_array;
  assign w_array = {prot_w,T_432};
  assign T_433 = priv_ok & sx_array;
  assign x_array = {prot_x,T_433};
  assign T_435 = io_ptw_status_mxr ? xr_array : 4'h0;
  assign T_436 = sr_array | T_435;
  assign T_437 = priv_ok & T_436;
  assign r_array = {prot_r,T_437};
  assign c_array = {T_261,cash_array};
  assign T_438 = io_req_bits_vpn[27];
  assign T_439 = io_req_bits_vpn[26];
  assign bad_va = T_438 != T_439;
  assign T_467 = 2'h1 << 1'h1;
  assign GEN_32 = {{2'd0}, T_467};
  assign T_468 = T_403 | GEN_32;
  assign T_478 = 4'h1 << 2'h2;
  assign T_479 = T_468 | T_478;
  assign GEN_28 = io_req_valid ? T_479 : T_403;
  assign T_485 = state == 2'h0;
  assign T_486 = ~ r_array;
  assign T_487 = T_486 & 5'h10;
  assign T_489 = T_487 != 5'h0;
  assign T_490 = bad_va | T_489;
  assign T_491 = ~ w_array;
  assign T_492 = T_491 & 5'h10;
  assign T_494 = T_492 != 5'h0;
  assign T_495 = bad_va | T_494;
  assign T_496 = ~ x_array;
  assign T_497 = T_496 & 5'h10;
  assign T_499 = T_497 != 5'h0;
  assign T_500 = bad_va | T_499;
  assign T_501 = c_array & 5'h10;
  assign T_503 = T_501 != 5'h0;
  assign T_520 = passthrough_ppn;
  assign T_521 = state == 2'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  valid = GEN_2[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  ppns_0 = GEN_3[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {1{$random}};
  ppns_1 = GEN_4[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  ppns_2 = GEN_5[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  ppns_3 = GEN_6[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {2{$random}};
  tags_0 = GEN_7[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {2{$random}};
  tags_1 = GEN_8[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {2{$random}};
  tags_2 = GEN_9[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {2{$random}};
  tags_3 = GEN_10[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_11 = {1{$random}};
  state = GEN_11[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_12 = {2{$random}};
  r_refill_tag = GEN_12[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_13 = {1{$random}};
  r_refill_waddr = GEN_13[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_14 = {1{$random}};
  r_req_vpn = GEN_14[27:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_15 = {1{$random}};
  r_req_passthrough = GEN_15[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_16 = {1{$random}};
  r_req_instruction = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {1{$random}};
  r_req_store = GEN_17[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {1{$random}};
  pte_array_reserved_for_hardware = GEN_18[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_19 = {2{$random}};
  pte_array_ppn = GEN_19[37:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_20 = {1{$random}};
  pte_array_reserved_for_software = GEN_20[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_21 = {1{$random}};
  pte_array_d = GEN_21[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_22 = {1{$random}};
  pte_array_a = GEN_22[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_23 = {1{$random}};
  pte_array_g = GEN_23[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_24 = {1{$random}};
  pte_array_u = GEN_24[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_25 = {1{$random}};
  pte_array_x = GEN_25[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_26 = {1{$random}};
  pte_array_w = GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_27 = {1{$random}};
  pte_array_r = GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  pte_array_v = GEN_30[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  u_array = GEN_31[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  sw_array = GEN_33[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  sx_array = GEN_34[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {1{$random}};
  sr_array = GEN_35[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  xr_array = GEN_36[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  cash_array = GEN_37[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {1{$random}};
  dirty_array = GEN_38[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  T_403 = GEN_39[3:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      valid <= 4'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(reset) begin
      state <= 2'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(io_req_valid) begin
        T_403 <= T_479;
      end
    end
  end
endmodule
module Frontend(
  input   clk,
  input   reset,
  input   io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_pc,
  input   io_cpu_req_bits_speculative,
  input   io_cpu_resp_ready,
  output  io_cpu_resp_valid,
  output  io_cpu_resp_bits_btb_valid,
  output  io_cpu_resp_bits_btb_bits_taken,
  output [1:0] io_cpu_resp_bits_btb_bits_mask,
  output  io_cpu_resp_bits_btb_bits_bridx,
  output [38:0] io_cpu_resp_bits_btb_bits_target,
  output  io_cpu_resp_bits_btb_bits_entry,
  output  io_cpu_resp_bits_btb_bits_bht_history,
  output [1:0] io_cpu_resp_bits_btb_bits_bht_value,
  output [39:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data,
  output [1:0] io_cpu_resp_bits_mask,
  output  io_cpu_resp_bits_xcpt_if,
  output  io_cpu_resp_bits_replay,
  input   io_cpu_btb_update_valid,
  input   io_cpu_btb_update_bits_prediction_valid,
  input   io_cpu_btb_update_bits_prediction_bits_taken,
  input  [1:0] io_cpu_btb_update_bits_prediction_bits_mask,
  input   io_cpu_btb_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_btb_update_bits_prediction_bits_target,
  input   io_cpu_btb_update_bits_prediction_bits_entry,
  input   io_cpu_btb_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
  input  [38:0] io_cpu_btb_update_bits_pc,
  input  [38:0] io_cpu_btb_update_bits_target,
  input   io_cpu_btb_update_bits_taken,
  input   io_cpu_btb_update_bits_isValid,
  input   io_cpu_btb_update_bits_isJump,
  input   io_cpu_btb_update_bits_isReturn,
  input  [38:0] io_cpu_btb_update_bits_br_pc,
  input   io_cpu_bht_update_valid,
  input   io_cpu_bht_update_bits_prediction_valid,
  input   io_cpu_bht_update_bits_prediction_bits_taken,
  input  [1:0] io_cpu_bht_update_bits_prediction_bits_mask,
  input   io_cpu_bht_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_bht_update_bits_prediction_bits_target,
  input   io_cpu_bht_update_bits_prediction_bits_entry,
  input   io_cpu_bht_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
  input  [38:0] io_cpu_bht_update_bits_pc,
  input   io_cpu_bht_update_bits_taken,
  input   io_cpu_bht_update_bits_mispredict,
  input   io_cpu_ras_update_valid,
  input   io_cpu_ras_update_bits_isCall,
  input   io_cpu_ras_update_bits_isReturn,
  input  [38:0] io_cpu_ras_update_bits_returnAddr,
  input   io_cpu_ras_update_bits_prediction_valid,
  input   io_cpu_ras_update_bits_prediction_bits_taken,
  input  [1:0] io_cpu_ras_update_bits_prediction_bits_mask,
  input   io_cpu_ras_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_ras_update_bits_prediction_bits_target,
  input   io_cpu_ras_update_bits_prediction_bits_entry,
  input   io_cpu_ras_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
  input   io_cpu_flush_icache,
  input   io_cpu_flush_tlb,
  output [39:0] io_cpu_npc,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_pum,
  output  io_ptw_req_bits_mxr,
  output [26:0] io_ptw_req_bits_addr,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [15:0] io_ptw_resp_bits_pte_reserved_for_hardware,
  input  [37:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_a,
  input   io_ptw_resp_bits_pte_g,
  input   io_ptw_resp_bits_pte_u,
  input   io_ptw_resp_bits_pte_x,
  input   io_ptw_resp_bits_pte_w,
  input   io_ptw_resp_bits_pte_r,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [37:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [3:0] io_ptw_status_zero1,
  input   io_ptw_status_mxr,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output  io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [10:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input   io_mem_grant_bits_client_xact_id,
  input  [1:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_req_valid;
  wire [38:0] icache_io_req_bits_addr;
  wire [19:0] icache_io_s1_ppn;
  wire  icache_io_s1_kill;
  wire  icache_io_s2_kill;
  wire  icache_io_resp_ready;
  wire  icache_io_resp_valid;
  wire [15:0] icache_io_resp_bits_data;
  wire [63:0] icache_io_resp_bits_datablock;
  wire  icache_io_invalidate;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire  icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [10:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire  icache_io_mem_grant_bits_client_xact_id;
  wire [1:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  tlb_clk;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [27:0] tlb_io_req_bits_vpn;
  wire  tlb_io_req_bits_passthrough;
  wire  tlb_io_req_bits_instruction;
  wire  tlb_io_req_bits_store;
  wire  tlb_io_resp_miss;
  wire [19:0] tlb_io_resp_ppn;
  wire  tlb_io_resp_xcpt_ld;
  wire  tlb_io_resp_xcpt_st;
  wire  tlb_io_resp_xcpt_if;
  wire  tlb_io_resp_cacheable;
  wire  tlb_io_ptw_req_ready;
  wire  tlb_io_ptw_req_valid;
  wire [1:0] tlb_io_ptw_req_bits_prv;
  wire  tlb_io_ptw_req_bits_pum;
  wire  tlb_io_ptw_req_bits_mxr;
  wire [26:0] tlb_io_ptw_req_bits_addr;
  wire  tlb_io_ptw_req_bits_store;
  wire  tlb_io_ptw_req_bits_fetch;
  wire  tlb_io_ptw_resp_valid;
  wire [15:0] tlb_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] tlb_io_ptw_resp_bits_pte_ppn;
  wire [1:0] tlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  tlb_io_ptw_resp_bits_pte_d;
  wire  tlb_io_ptw_resp_bits_pte_a;
  wire  tlb_io_ptw_resp_bits_pte_g;
  wire  tlb_io_ptw_resp_bits_pte_u;
  wire  tlb_io_ptw_resp_bits_pte_x;
  wire  tlb_io_ptw_resp_bits_pte_w;
  wire  tlb_io_ptw_resp_bits_pte_r;
  wire  tlb_io_ptw_resp_bits_pte_v;
  wire [6:0] tlb_io_ptw_ptbr_asid;
  wire [37:0] tlb_io_ptw_ptbr_ppn;
  wire  tlb_io_ptw_invalidate;
  wire  tlb_io_ptw_status_debug;
  wire [1:0] tlb_io_ptw_status_prv;
  wire  tlb_io_ptw_status_sd;
  wire [30:0] tlb_io_ptw_status_zero3;
  wire  tlb_io_ptw_status_sd_rv32;
  wire [1:0] tlb_io_ptw_status_zero2;
  wire [4:0] tlb_io_ptw_status_vm;
  wire [3:0] tlb_io_ptw_status_zero1;
  wire  tlb_io_ptw_status_mxr;
  wire  tlb_io_ptw_status_pum;
  wire  tlb_io_ptw_status_mprv;
  wire [1:0] tlb_io_ptw_status_xs;
  wire [1:0] tlb_io_ptw_status_fs;
  wire [1:0] tlb_io_ptw_status_mpp;
  wire [1:0] tlb_io_ptw_status_hpp;
  wire  tlb_io_ptw_status_spp;
  wire  tlb_io_ptw_status_mpie;
  wire  tlb_io_ptw_status_hpie;
  wire  tlb_io_ptw_status_spie;
  wire  tlb_io_ptw_status_upie;
  wire  tlb_io_ptw_status_mie;
  wire  tlb_io_ptw_status_hie;
  wire  tlb_io_ptw_status_sie;
  wire  tlb_io_ptw_status_uie;
  reg [39:0] s1_pc_;
  reg [63:0] GEN_17;
  wire [39:0] T_1483;
  wire [39:0] T_1485;
  wire [39:0] s1_pc;
  reg  s1_speculative;
  reg [31:0] GEN_18;
  reg  s1_same_block;
  reg [31:0] GEN_19;
  reg  s2_valid;
  reg [31:0] GEN_20;
  reg [39:0] s2_pc;
  reg [63:0] GEN_21;
  reg  s2_btb_resp_valid;
  reg [31:0] GEN_22;
  reg  s2_btb_resp_bits_taken;
  reg [31:0] GEN_23;
  reg [1:0] s2_btb_resp_bits_mask;
  reg [31:0] GEN_24;
  reg  s2_btb_resp_bits_bridx;
  reg [31:0] GEN_25;
  reg [38:0] s2_btb_resp_bits_target;
  reg [63:0] GEN_26;
  reg  s2_btb_resp_bits_entry;
  reg [31:0] GEN_27;
  reg  s2_btb_resp_bits_bht_history;
  reg [31:0] GEN_28;
  reg [1:0] s2_btb_resp_bits_bht_value;
  reg [31:0] GEN_29;
  reg  s2_xcpt_if;
  reg [31:0] GEN_30;
  reg  s2_speculative;
  reg [31:0] GEN_31;
  reg  s2_cacheable;
  reg [31:0] GEN_32;
  wire [39:0] T_1511;
  wire [39:0] T_1513;
  wire [39:0] T_1514;
  wire [40:0] T_1516;
  wire [39:0] ntpc;
  wire [39:0] T_1518;
  wire [39:0] T_1520;
  wire  ntpc_same_block;
  wire [39:0] predicted_npc;
  wire  predicted_taken;
  wire  T_1523;
  wire  icmiss;
  wire [39:0] npc;
  wire  T_1525;
  wire  T_1527;
  wire  T_1528;
  wire  T_1530;
  wire  T_1531;
  wire  s0_same_block;
  wire  T_1533;
  wire  stall;
  wire  T_1535;
  wire  T_1537;
  wire  T_1538;
  wire  T_1540;
  wire  T_1541;
  wire  T_1542;
  wire  T_1543;
  wire  T_1544;
  wire [39:0] GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire [39:0] GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [39:0] GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [39:0] GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  T_1555;
  wire [27:0] T_1556;
  wire  T_1563;
  wire  T_1564;
  wire  T_1565;
  wire  T_1566;
  wire  T_1567;
  wire  T_1568;
  wire  T_1570;
  wire  T_1571;
  wire  T_1575;
  wire  T_1576;
  wire  T_1577;
  wire  T_1578;
  wire  T_1579;
  wire [39:0] T_1580;
  wire  T_1581;
  wire [5:0] GEN_16;
  wire [5:0] T_1582;
  wire [63:0] T_1583;
  wire  T_1585;
  wire [2:0] T_1586;
  wire  T_1589;
  wire  T_1591;
  wire  T_1592;
  ICache icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_ppn(icache_io_s1_ppn),
    .io_s1_kill(icache_io_s1_kill),
    .io_s2_kill(icache_io_s2_kill),
    .io_resp_ready(icache_io_resp_ready),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_datablock(icache_io_resp_bits_datablock),
    .io_invalidate(icache_io_invalidate),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  TLB tlb (
    .clk(tlb_clk),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vpn(tlb_io_req_bits_vpn),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_instruction(tlb_io_req_bits_instruction),
    .io_req_bits_store(tlb_io_req_bits_store),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_ppn(tlb_io_resp_ppn),
    .io_resp_xcpt_ld(tlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(tlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(tlb_io_resp_xcpt_if),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_prv(tlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(tlb_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(tlb_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(tlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(tlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(tlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(tlb_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(tlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(tlb_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(tlb_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(tlb_io_ptw_invalidate),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_status_sd(tlb_io_ptw_status_sd),
    .io_ptw_status_zero3(tlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(tlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(tlb_io_ptw_status_zero2),
    .io_ptw_status_vm(tlb_io_ptw_status_vm),
    .io_ptw_status_zero1(tlb_io_ptw_status_zero1),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_pum(tlb_io_ptw_status_pum),
    .io_ptw_status_mprv(tlb_io_ptw_status_mprv),
    .io_ptw_status_xs(tlb_io_ptw_status_xs),
    .io_ptw_status_fs(tlb_io_ptw_status_fs),
    .io_ptw_status_mpp(tlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(tlb_io_ptw_status_hpp),
    .io_ptw_status_spp(tlb_io_ptw_status_spp),
    .io_ptw_status_mpie(tlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(tlb_io_ptw_status_hpie),
    .io_ptw_status_spie(tlb_io_ptw_status_spie),
    .io_ptw_status_upie(tlb_io_ptw_status_upie),
    .io_ptw_status_mie(tlb_io_ptw_status_mie),
    .io_ptw_status_hie(tlb_io_ptw_status_hie),
    .io_ptw_status_sie(tlb_io_ptw_status_sie),
    .io_ptw_status_uie(tlb_io_ptw_status_uie)
  );
  assign io_cpu_resp_valid = T_1579;
  assign io_cpu_resp_bits_btb_valid = s2_btb_resp_valid;
  assign io_cpu_resp_bits_btb_bits_taken = s2_btb_resp_bits_taken;
  assign io_cpu_resp_bits_btb_bits_mask = s2_btb_resp_bits_mask;
  assign io_cpu_resp_bits_btb_bits_bridx = s2_btb_resp_bits_bridx;
  assign io_cpu_resp_bits_btb_bits_target = s2_btb_resp_bits_target;
  assign io_cpu_resp_bits_btb_bits_entry = s2_btb_resp_bits_entry;
  assign io_cpu_resp_bits_btb_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign io_cpu_resp_bits_btb_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign io_cpu_resp_bits_pc = s2_pc;
  assign io_cpu_resp_bits_data = T_1583[31:0];
  assign io_cpu_resp_bits_mask = T_1586[1:0];
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign io_cpu_resp_bits_replay = T_1592;
  assign io_cpu_npc = T_1580;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_pum = tlb_io_ptw_req_bits_pum;
  assign io_ptw_req_bits_mxr = tlb_io_ptw_req_bits_mxr;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_mem_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_mem_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_mem_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_mem_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_mem_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_req_valid = T_1564;
  assign icache_io_req_bits_addr = io_cpu_npc[38:0];
  assign icache_io_s1_ppn = tlb_io_resp_ppn;
  assign icache_io_s1_kill = T_1568;
  assign icache_io_s2_kill = T_1571;
  assign icache_io_resp_ready = T_1576;
  assign icache_io_invalidate = io_cpu_flush_icache;
  assign icache_io_mem_acquire_ready = io_mem_acquire_ready;
  assign icache_io_mem_grant_valid = io_mem_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign tlb_clk = clk;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = T_1555;
  assign tlb_io_req_bits_vpn = T_1556;
  assign tlb_io_req_bits_passthrough = 1'h0;
  assign tlb_io_req_bits_instruction = 1'h1;
  assign tlb_io_req_bits_store = 1'h0;
  assign tlb_io_ptw_req_ready = io_ptw_req_ready;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_hardware = io_ptw_resp_bits_pte_reserved_for_hardware;
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a;
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g;
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u;
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x;
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w;
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign tlb_io_ptw_ptbr_asid = io_ptw_ptbr_asid;
  assign tlb_io_ptw_ptbr_ppn = io_ptw_ptbr_ppn;
  assign tlb_io_ptw_invalidate = io_ptw_invalidate;
  assign tlb_io_ptw_status_debug = io_ptw_status_debug;
  assign tlb_io_ptw_status_prv = io_ptw_status_prv;
  assign tlb_io_ptw_status_sd = io_ptw_status_sd;
  assign tlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign tlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign tlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign tlb_io_ptw_status_vm = io_ptw_status_vm;
  assign tlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr;
  assign tlb_io_ptw_status_pum = io_ptw_status_pum;
  assign tlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign tlb_io_ptw_status_xs = io_ptw_status_xs;
  assign tlb_io_ptw_status_fs = io_ptw_status_fs;
  assign tlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign tlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign tlb_io_ptw_status_spp = io_ptw_status_spp;
  assign tlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign tlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign tlb_io_ptw_status_spie = io_ptw_status_spie;
  assign tlb_io_ptw_status_upie = io_ptw_status_upie;
  assign tlb_io_ptw_status_mie = io_ptw_status_mie;
  assign tlb_io_ptw_status_hie = io_ptw_status_hie;
  assign tlb_io_ptw_status_sie = io_ptw_status_sie;
  assign tlb_io_ptw_status_uie = io_ptw_status_uie;
  assign T_1483 = ~ s1_pc_;
  assign T_1485 = T_1483 | 40'h1;
  assign s1_pc = ~ T_1485;
  assign T_1511 = ~ s1_pc;
  assign T_1513 = T_1511 | 40'h3;
  assign T_1514 = ~ T_1513;
  assign T_1516 = T_1514 + 40'h4;
  assign ntpc = T_1516[39:0];
  assign T_1518 = ntpc & 40'h8;
  assign T_1520 = s1_pc & 40'h8;
  assign ntpc_same_block = T_1518 == T_1520;
  assign predicted_npc = ntpc;
  assign predicted_taken = 1'h0;
  assign T_1523 = icache_io_resp_valid == 1'h0;
  assign icmiss = s2_valid & T_1523;
  assign npc = icmiss ? s2_pc : predicted_npc;
  assign T_1525 = predicted_taken == 1'h0;
  assign T_1527 = icmiss == 1'h0;
  assign T_1528 = T_1525 & T_1527;
  assign T_1530 = io_cpu_req_valid == 1'h0;
  assign T_1531 = T_1528 & T_1530;
  assign s0_same_block = T_1531 & ntpc_same_block;
  assign T_1533 = io_cpu_resp_ready == 1'h0;
  assign stall = io_cpu_resp_valid & T_1533;
  assign T_1535 = stall == 1'h0;
  assign T_1537 = tlb_io_resp_miss == 1'h0;
  assign T_1538 = s0_same_block & T_1537;
  assign T_1540 = s2_speculative == 1'h0;
  assign T_1541 = s2_valid & T_1540;
  assign T_1542 = s1_speculative | T_1541;
  assign T_1543 = T_1542 | predicted_taken;
  assign T_1544 = icmiss ? s2_speculative : T_1543;
  assign GEN_0 = T_1527 ? s1_pc : s2_pc;
  assign GEN_1 = T_1527 ? s1_speculative : s2_speculative;
  assign GEN_2 = T_1527 ? tlb_io_resp_cacheable : s2_cacheable;
  assign GEN_3 = T_1527 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign GEN_4 = T_1535 ? T_1538 : s1_same_block;
  assign GEN_5 = T_1535 ? io_cpu_npc : s1_pc_;
  assign GEN_6 = T_1535 ? T_1544 : s1_speculative;
  assign GEN_7 = T_1535 ? T_1527 : s2_valid;
  assign GEN_8 = T_1535 ? GEN_0 : s2_pc;
  assign GEN_9 = T_1535 ? GEN_1 : s2_speculative;
  assign GEN_10 = T_1535 ? GEN_2 : s2_cacheable;
  assign GEN_11 = T_1535 ? GEN_3 : s2_xcpt_if;
  assign GEN_12 = io_cpu_req_valid ? 1'h0 : GEN_4;
  assign GEN_13 = io_cpu_req_valid ? io_cpu_npc : GEN_5;
  assign GEN_14 = io_cpu_req_valid ? io_cpu_req_bits_speculative : GEN_6;
  assign GEN_15 = io_cpu_req_valid ? 1'h0 : GEN_7;
  assign T_1555 = T_1535 & T_1527;
  assign T_1556 = s1_pc[39:12];
  assign T_1563 = s0_same_block == 1'h0;
  assign T_1564 = T_1535 & T_1563;
  assign T_1565 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T_1566 = T_1565 | tlb_io_resp_xcpt_if;
  assign T_1567 = T_1566 | icmiss;
  assign T_1568 = T_1567 | io_cpu_flush_tlb;
  assign T_1570 = s2_cacheable == 1'h0;
  assign T_1571 = s2_speculative & T_1570;
  assign T_1575 = s1_same_block == 1'h0;
  assign T_1576 = T_1535 & T_1575;
  assign T_1577 = icache_io_resp_valid | icache_io_s2_kill;
  assign T_1578 = T_1577 | s2_xcpt_if;
  assign T_1579 = s2_valid & T_1578;
  assign T_1580 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign T_1581 = s2_pc[2];
  assign GEN_16 = {{5'd0}, T_1581};
  assign T_1582 = GEN_16 << 5;
  assign T_1583 = icache_io_resp_bits_datablock >> T_1582;
  assign T_1585 = s2_pc[1];
  assign T_1586 = 3'h3 << T_1585;
  assign T_1589 = icache_io_s2_kill & T_1523;
  assign T_1591 = s2_xcpt_if == 1'h0;
  assign T_1592 = T_1589 & T_1591;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {2{$random}};
  s1_pc_ = GEN_17[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {1{$random}};
  s1_speculative = GEN_18[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_19 = {1{$random}};
  s1_same_block = GEN_19[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_20 = {1{$random}};
  s2_valid = GEN_20[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_21 = {2{$random}};
  s2_pc = GEN_21[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_22 = {1{$random}};
  s2_btb_resp_valid = GEN_22[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_23 = {1{$random}};
  s2_btb_resp_bits_taken = GEN_23[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_24 = {1{$random}};
  s2_btb_resp_bits_mask = GEN_24[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_25 = {1{$random}};
  s2_btb_resp_bits_bridx = GEN_25[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_26 = {2{$random}};
  s2_btb_resp_bits_target = GEN_26[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_27 = {1{$random}};
  s2_btb_resp_bits_entry = GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_28 = {1{$random}};
  s2_btb_resp_bits_bht_history = GEN_28[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  s2_btb_resp_bits_bht_value = GEN_29[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  s2_xcpt_if = GEN_30[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  s2_speculative = GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  s2_cacheable = GEN_32[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_pc_ <= io_cpu_npc;
      end else begin
        if(T_1535) begin
          s1_pc_ <= io_cpu_npc;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_speculative <= io_cpu_req_bits_speculative;
      end else begin
        if(T_1535) begin
          if(icmiss) begin
            s1_speculative <= s2_speculative;
          end else begin
            s1_speculative <= T_1543;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_same_block <= 1'h0;
      end else begin
        if(T_1535) begin
          s1_same_block <= T_1538;
        end
      end
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else begin
      if(io_cpu_req_valid) begin
        s2_valid <= 1'h0;
      end else begin
        if(T_1535) begin
          s2_valid <= T_1527;
        end
      end
    end
    if(reset) begin
      s2_pc <= 40'h1000;
    end else begin
      if(T_1535) begin
        if(T_1527) begin
          s2_pc <= s1_pc;
        end
      end
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else begin
      if(T_1535) begin
        if(T_1527) begin
          s2_xcpt_if <= tlb_io_resp_xcpt_if;
        end
      end
    end
    if(reset) begin
      s2_speculative <= 1'h0;
    end else begin
      if(T_1535) begin
        if(T_1527) begin
          s2_speculative <= s1_speculative;
        end
      end
    end
    if(reset) begin
      s2_cacheable <= 1'h0;
    end else begin
      if(T_1535) begin
        if(T_1527) begin
          s2_cacheable <= tlb_io_resp_cacheable;
        end
      end
    end
  end
endmodule
module FinishQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output  io_count
);
  reg [1:0] ram_manager_xact_id [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_manager_xact_id_T_254_data;
  wire  ram_manager_xact_id_T_254_addr;
  wire  ram_manager_xact_id_T_254_en;
  wire [1:0] ram_manager_xact_id_T_224_data;
  wire  ram_manager_xact_id_T_224_addr;
  wire  ram_manager_xact_id_T_224_mask;
  wire  ram_manager_xact_id_T_224_en;
  reg  ram_manager_id [0:0];
  reg [31:0] GEN_1;
  wire  ram_manager_id_T_254_data;
  wire  ram_manager_id_T_254_addr;
  wire  ram_manager_id_T_254_en;
  wire  ram_manager_id_T_224_data;
  wire  ram_manager_id_T_224_addr;
  wire  ram_manager_id_T_224_mask;
  wire  ram_manager_id_T_224_en;
  reg  maybe_full;
  reg [31:0] GEN_2;
  wire  T_221;
  wire  T_222;
  wire  do_enq;
  wire  T_223;
  wire  do_deq;
  wire  T_249;
  wire  GEN_7;
  wire  T_251;
  wire [1:0] T_277;
  wire  ptr_diff;
  wire [1:0] T_279;
  assign io_enq_ready = T_221;
  assign io_deq_valid = T_251;
  assign io_deq_bits_manager_xact_id = ram_manager_xact_id_T_254_data;
  assign io_deq_bits_manager_id = ram_manager_id_T_254_data;
  assign io_count = T_279[0];
  assign ram_manager_xact_id_T_254_addr = 1'h0;
  assign ram_manager_xact_id_T_254_en = 1'h1;
  assign ram_manager_xact_id_T_254_data = ram_manager_xact_id[ram_manager_xact_id_T_254_addr];
  assign ram_manager_xact_id_T_224_data = io_enq_bits_manager_xact_id;
  assign ram_manager_xact_id_T_224_addr = 1'h0;
  assign ram_manager_xact_id_T_224_mask = do_enq;
  assign ram_manager_xact_id_T_224_en = do_enq;
  assign ram_manager_id_T_254_addr = 1'h0;
  assign ram_manager_id_T_254_en = 1'h1;
  assign ram_manager_id_T_254_data = ram_manager_id[ram_manager_id_T_254_addr];
  assign ram_manager_id_T_224_data = io_enq_bits_manager_id;
  assign ram_manager_id_T_224_addr = 1'h0;
  assign ram_manager_id_T_224_mask = do_enq;
  assign ram_manager_id_T_224_en = do_enq;
  assign T_221 = maybe_full == 1'h0;
  assign T_222 = io_enq_ready & io_enq_valid;
  assign do_enq = T_222;
  assign T_223 = io_deq_ready & io_deq_valid;
  assign do_deq = T_223;
  assign T_249 = do_enq != do_deq;
  assign GEN_7 = T_249 ? do_enq : maybe_full;
  assign T_251 = T_221 == 1'h0;
  assign T_277 = 1'h0 - 1'h0;
  assign ptr_diff = T_277[0:0];
  assign T_279 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_manager_xact_id[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_manager_id[initvar] = GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  maybe_full = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_manager_xact_id_T_224_en & ram_manager_xact_id_T_224_mask) begin
      ram_manager_xact_id[ram_manager_xact_id_T_224_addr] <= ram_manager_xact_id_T_224_data;
    end
    if(ram_manager_id_T_224_en & ram_manager_id_T_224_mask) begin
      ram_manager_id[ram_manager_id_T_224_addr] <= ram_manager_id_T_224_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_249) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Arbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input   io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input   io_in_1_bits_way_en,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [5:0] io_in_2_bits_idx,
  input   io_in_2_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output  io_out_bits_way_en,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [5:0] GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [5:0] GEN_4;
  wire  GEN_5;
  wire  T_637;
  wire  grant_1;
  wire  grant_2;
  wire  T_641;
  wire  T_642;
  wire  T_644;
  wire  T_645;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_641;
  assign io_in_2_ready = T_642;
  assign io_out_valid = T_645;
  assign io_out_bits_idx = GEN_4;
  assign io_out_bits_way_en = GEN_5;
  assign io_chosen = GEN_3;
  assign GEN_0 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_1 = io_in_1_valid ? io_in_1_bits_idx : io_in_2_bits_idx;
  assign GEN_2 = io_in_1_valid ? io_in_1_bits_way_en : io_in_2_bits_way_en;
  assign GEN_3 = io_in_0_valid ? 2'h0 : GEN_0;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_idx : GEN_1;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_way_en : GEN_2;
  assign T_637 = io_in_0_valid | io_in_1_valid;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign grant_2 = T_637 == 1'h0;
  assign T_641 = grant_1 & io_out_ready;
  assign T_642 = grant_2 & io_out_ready;
  assign T_644 = grant_2 == 1'h0;
  assign T_645 = T_644 | io_in_2_valid;
endmodule
module Arbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input   io_in_0_bits_way_en,
  input  [19:0] io_in_0_bits_data_tag,
  input  [1:0] io_in_0_bits_data_coh_state,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input   io_in_1_bits_way_en,
  input  [19:0] io_in_1_bits_data_tag,
  input  [1:0] io_in_1_bits_data_coh_state,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [5:0] io_in_2_bits_idx,
  input   io_in_2_bits_way_en,
  input  [19:0] io_in_2_bits_data_tag,
  input  [1:0] io_in_2_bits_data_coh_state,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output  io_out_bits_way_en,
  output [19:0] io_out_bits_data_tag,
  output [1:0] io_out_bits_data_coh_state,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [5:0] GEN_1;
  wire  GEN_2;
  wire [19:0] GEN_3;
  wire [1:0] GEN_4;
  wire [1:0] GEN_5;
  wire [5:0] GEN_6;
  wire  GEN_7;
  wire [19:0] GEN_8;
  wire [1:0] GEN_9;
  wire  T_2821;
  wire  grant_1;
  wire  grant_2;
  wire  T_2825;
  wire  T_2826;
  wire  T_2828;
  wire  T_2829;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_2825;
  assign io_in_2_ready = T_2826;
  assign io_out_valid = T_2829;
  assign io_out_bits_idx = GEN_6;
  assign io_out_bits_way_en = GEN_7;
  assign io_out_bits_data_tag = GEN_8;
  assign io_out_bits_data_coh_state = GEN_9;
  assign io_chosen = GEN_5;
  assign GEN_0 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_1 = io_in_1_valid ? io_in_1_bits_idx : io_in_2_bits_idx;
  assign GEN_2 = io_in_1_valid ? io_in_1_bits_way_en : io_in_2_bits_way_en;
  assign GEN_3 = io_in_1_valid ? io_in_1_bits_data_tag : io_in_2_bits_data_tag;
  assign GEN_4 = io_in_1_valid ? io_in_1_bits_data_coh_state : io_in_2_bits_data_coh_state;
  assign GEN_5 = io_in_0_valid ? 2'h0 : GEN_0;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_idx : GEN_1;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_way_en : GEN_2;
  assign GEN_8 = io_in_0_valid ? io_in_0_bits_data_tag : GEN_3;
  assign GEN_9 = io_in_0_valid ? io_in_0_bits_data_coh_state : GEN_4;
  assign T_2821 = io_in_0_valid | io_in_1_valid;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign grant_2 = T_2821 == 1'h0;
  assign T_2825 = grant_1 & io_out_ready;
  assign T_2826 = grant_2 & io_out_ready;
  assign T_2828 = grant_2 == 1'h0;
  assign T_2829 = T_2828 | io_in_2_valid;
endmodule
module DCacheDataArray(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [11:0] io_req_bits_addr,
  input   io_req_bits_write,
  input  [63:0] io_req_bits_wdata,
  input  [7:0] io_req_bits_wmask,
  input   io_req_bits_way_en,
  output [63:0] io_resp_0
);
  wire [8:0] addr;
  reg [7:0] T_406_0 [0:511];
  reg [31:0] GEN_0;
  wire [7:0] T_406_0_T_446_data;
  wire [8:0] T_406_0_T_446_addr;
  wire  T_406_0_T_446_en;
  reg [8:0] GEN_1;
  reg [31:0] GEN_2;
  wire [7:0] T_406_0_T_437_data;
  wire [8:0] T_406_0_T_437_addr;
  wire  T_406_0_T_437_mask;
  wire  T_406_0_T_437_en;
  reg [7:0] T_406_1 [0:511];
  reg [31:0] GEN_3;
  wire [7:0] T_406_1_T_446_data;
  wire [8:0] T_406_1_T_446_addr;
  wire  T_406_1_T_446_en;
  reg [8:0] GEN_4;
  reg [31:0] GEN_5;
  wire [7:0] T_406_1_T_437_data;
  wire [8:0] T_406_1_T_437_addr;
  wire  T_406_1_T_437_mask;
  wire  T_406_1_T_437_en;
  reg [7:0] T_406_2 [0:511];
  reg [31:0] GEN_6;
  wire [7:0] T_406_2_T_446_data;
  wire [8:0] T_406_2_T_446_addr;
  wire  T_406_2_T_446_en;
  reg [8:0] GEN_7;
  reg [31:0] GEN_8;
  wire [7:0] T_406_2_T_437_data;
  wire [8:0] T_406_2_T_437_addr;
  wire  T_406_2_T_437_mask;
  wire  T_406_2_T_437_en;
  reg [7:0] T_406_3 [0:511];
  reg [31:0] GEN_9;
  wire [7:0] T_406_3_T_446_data;
  wire [8:0] T_406_3_T_446_addr;
  wire  T_406_3_T_446_en;
  reg [8:0] GEN_10;
  reg [31:0] GEN_11;
  wire [7:0] T_406_3_T_437_data;
  wire [8:0] T_406_3_T_437_addr;
  wire  T_406_3_T_437_mask;
  wire  T_406_3_T_437_en;
  reg [7:0] T_406_4 [0:511];
  reg [31:0] GEN_12;
  wire [7:0] T_406_4_T_446_data;
  wire [8:0] T_406_4_T_446_addr;
  wire  T_406_4_T_446_en;
  reg [8:0] GEN_13;
  reg [31:0] GEN_14;
  wire [7:0] T_406_4_T_437_data;
  wire [8:0] T_406_4_T_437_addr;
  wire  T_406_4_T_437_mask;
  wire  T_406_4_T_437_en;
  reg [7:0] T_406_5 [0:511];
  reg [31:0] GEN_15;
  wire [7:0] T_406_5_T_446_data;
  wire [8:0] T_406_5_T_446_addr;
  wire  T_406_5_T_446_en;
  reg [8:0] GEN_16;
  reg [31:0] GEN_17;
  wire [7:0] T_406_5_T_437_data;
  wire [8:0] T_406_5_T_437_addr;
  wire  T_406_5_T_437_mask;
  wire  T_406_5_T_437_en;
  reg [7:0] T_406_6 [0:511];
  reg [31:0] GEN_18;
  wire [7:0] T_406_6_T_446_data;
  wire [8:0] T_406_6_T_446_addr;
  wire  T_406_6_T_446_en;
  reg [8:0] GEN_19;
  reg [31:0] GEN_20;
  wire [7:0] T_406_6_T_437_data;
  wire [8:0] T_406_6_T_437_addr;
  wire  T_406_6_T_437_mask;
  wire  T_406_6_T_437_en;
  reg [7:0] T_406_7 [0:511];
  reg [31:0] GEN_21;
  wire [7:0] T_406_7_T_446_data;
  wire [8:0] T_406_7_T_446_addr;
  wire  T_406_7_T_446_en;
  reg [8:0] GEN_22;
  reg [31:0] GEN_23;
  wire [7:0] T_406_7_T_437_data;
  wire [8:0] T_406_7_T_437_addr;
  wire  T_406_7_T_437_mask;
  wire  T_406_7_T_437_en;
  wire  T_411;
  wire [7:0] T_412;
  wire [7:0] T_413;
  wire [7:0] T_414;
  wire [7:0] T_415;
  wire [7:0] T_416;
  wire [7:0] T_417;
  wire [7:0] T_418;
  wire [7:0] T_419;
  wire [7:0] T_425_0;
  wire [7:0] T_425_1;
  wire [7:0] T_425_2;
  wire [7:0] T_425_3;
  wire [7:0] T_425_4;
  wire [7:0] T_425_5;
  wire [7:0] T_425_6;
  wire [7:0] T_425_7;
  wire  T_427;
  wire  T_428;
  wire  T_429;
  wire  T_430;
  wire  T_431;
  wire  T_432;
  wire  T_433;
  wire  T_434;
  wire  GEN_28;
  wire  GEN_30;
  wire  GEN_32;
  wire  GEN_34;
  wire  GEN_36;
  wire  GEN_38;
  wire  GEN_40;
  wire  GEN_42;
  wire  T_440;
  wire  T_441;
  wire [8:0] T_443;
  wire [15:0] T_448;
  wire [15:0] T_449;
  wire [31:0] T_450;
  wire [15:0] T_451;
  wire [15:0] T_452;
  wire [31:0] T_453;
  wire [63:0] T_454;
  assign io_resp_0 = T_454;
  assign addr = io_req_bits_addr[11:3];
  assign T_406_0_T_446_addr = T_443;
  assign T_406_0_T_446_en = T_441;
  assign T_406_0_T_446_data = T_406_0[GEN_1];
  assign T_406_0_T_437_data = T_425_0;
  assign T_406_0_T_437_addr = addr;
  assign T_406_0_T_437_mask = GEN_28;
  assign T_406_0_T_437_en = T_411;
  assign T_406_1_T_446_addr = T_443;
  assign T_406_1_T_446_en = T_441;
  assign T_406_1_T_446_data = T_406_1[GEN_4];
  assign T_406_1_T_437_data = T_425_1;
  assign T_406_1_T_437_addr = addr;
  assign T_406_1_T_437_mask = GEN_30;
  assign T_406_1_T_437_en = T_411;
  assign T_406_2_T_446_addr = T_443;
  assign T_406_2_T_446_en = T_441;
  assign T_406_2_T_446_data = T_406_2[GEN_7];
  assign T_406_2_T_437_data = T_425_2;
  assign T_406_2_T_437_addr = addr;
  assign T_406_2_T_437_mask = GEN_32;
  assign T_406_2_T_437_en = T_411;
  assign T_406_3_T_446_addr = T_443;
  assign T_406_3_T_446_en = T_441;
  assign T_406_3_T_446_data = T_406_3[GEN_10];
  assign T_406_3_T_437_data = T_425_3;
  assign T_406_3_T_437_addr = addr;
  assign T_406_3_T_437_mask = GEN_34;
  assign T_406_3_T_437_en = T_411;
  assign T_406_4_T_446_addr = T_443;
  assign T_406_4_T_446_en = T_441;
  assign T_406_4_T_446_data = T_406_4[GEN_13];
  assign T_406_4_T_437_data = T_425_4;
  assign T_406_4_T_437_addr = addr;
  assign T_406_4_T_437_mask = GEN_36;
  assign T_406_4_T_437_en = T_411;
  assign T_406_5_T_446_addr = T_443;
  assign T_406_5_T_446_en = T_441;
  assign T_406_5_T_446_data = T_406_5[GEN_16];
  assign T_406_5_T_437_data = T_425_5;
  assign T_406_5_T_437_addr = addr;
  assign T_406_5_T_437_mask = GEN_38;
  assign T_406_5_T_437_en = T_411;
  assign T_406_6_T_446_addr = T_443;
  assign T_406_6_T_446_en = T_441;
  assign T_406_6_T_446_data = T_406_6[GEN_19];
  assign T_406_6_T_437_data = T_425_6;
  assign T_406_6_T_437_addr = addr;
  assign T_406_6_T_437_mask = GEN_40;
  assign T_406_6_T_437_en = T_411;
  assign T_406_7_T_446_addr = T_443;
  assign T_406_7_T_446_en = T_441;
  assign T_406_7_T_446_data = T_406_7[GEN_22];
  assign T_406_7_T_437_data = T_425_7;
  assign T_406_7_T_437_addr = addr;
  assign T_406_7_T_437_mask = GEN_42;
  assign T_406_7_T_437_en = T_411;
  assign T_411 = io_req_valid & io_req_bits_write;
  assign T_412 = io_req_bits_wdata[7:0];
  assign T_413 = io_req_bits_wdata[15:8];
  assign T_414 = io_req_bits_wdata[23:16];
  assign T_415 = io_req_bits_wdata[31:24];
  assign T_416 = io_req_bits_wdata[39:32];
  assign T_417 = io_req_bits_wdata[47:40];
  assign T_418 = io_req_bits_wdata[55:48];
  assign T_419 = io_req_bits_wdata[63:56];
  assign T_425_0 = T_412;
  assign T_425_1 = T_413;
  assign T_425_2 = T_414;
  assign T_425_3 = T_415;
  assign T_425_4 = T_416;
  assign T_425_5 = T_417;
  assign T_425_6 = T_418;
  assign T_425_7 = T_419;
  assign T_427 = io_req_bits_wmask[0];
  assign T_428 = io_req_bits_wmask[1];
  assign T_429 = io_req_bits_wmask[2];
  assign T_430 = io_req_bits_wmask[3];
  assign T_431 = io_req_bits_wmask[4];
  assign T_432 = io_req_bits_wmask[5];
  assign T_433 = io_req_bits_wmask[6];
  assign T_434 = io_req_bits_wmask[7];
  assign GEN_28 = T_411 ? T_427 : 1'h0;
  assign GEN_30 = T_411 ? T_428 : 1'h0;
  assign GEN_32 = T_411 ? T_429 : 1'h0;
  assign GEN_34 = T_411 ? T_430 : 1'h0;
  assign GEN_36 = T_411 ? T_431 : 1'h0;
  assign GEN_38 = T_411 ? T_432 : 1'h0;
  assign GEN_40 = T_411 ? T_433 : 1'h0;
  assign GEN_42 = T_411 ? T_434 : 1'h0;
  assign T_440 = io_req_bits_write == 1'h0;
  assign T_441 = io_req_valid & T_440;
  assign T_443 = addr;
  assign T_448 = {T_406_1_T_446_data,T_406_0_T_446_data};
  assign T_449 = {T_406_3_T_446_data,T_406_2_T_446_data};
  assign T_450 = {T_449,T_448};
  assign T_451 = {T_406_5_T_446_data,T_406_4_T_446_data};
  assign T_452 = {T_406_7_T_446_data,T_406_6_T_446_data};
  assign T_453 = {T_452,T_451};
  assign T_454 = {T_453,T_450};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_406_0[initvar] = GEN_0[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  GEN_1 = GEN_2[8:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_406_1[initvar] = GEN_3[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  GEN_4 = GEN_5[8:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_406_2[initvar] = GEN_6[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  GEN_7 = GEN_8[8:0];
  `endif
  GEN_9 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_406_3[initvar] = GEN_9[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_11 = {1{$random}};
  GEN_10 = GEN_11[8:0];
  `endif
  GEN_12 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_406_4[initvar] = GEN_12[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_14 = {1{$random}};
  GEN_13 = GEN_14[8:0];
  `endif
  GEN_15 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_406_5[initvar] = GEN_15[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {1{$random}};
  GEN_16 = GEN_17[8:0];
  `endif
  GEN_18 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_406_6[initvar] = GEN_18[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_20 = {1{$random}};
  GEN_19 = GEN_20[8:0];
  `endif
  GEN_21 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_406_7[initvar] = GEN_21[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_23 = {1{$random}};
  GEN_22 = GEN_23[8:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(T_406_0_T_446_en) begin
      GEN_1 <= T_406_0_T_446_addr;
    end
    if(T_406_0_T_437_en & T_406_0_T_437_mask) begin
      T_406_0[T_406_0_T_437_addr] <= T_406_0_T_437_data;
    end
    if(T_406_1_T_446_en) begin
      GEN_4 <= T_406_1_T_446_addr;
    end
    if(T_406_1_T_437_en & T_406_1_T_437_mask) begin
      T_406_1[T_406_1_T_437_addr] <= T_406_1_T_437_data;
    end
    if(T_406_2_T_446_en) begin
      GEN_7 <= T_406_2_T_446_addr;
    end
    if(T_406_2_T_437_en & T_406_2_T_437_mask) begin
      T_406_2[T_406_2_T_437_addr] <= T_406_2_T_437_data;
    end
    if(T_406_3_T_446_en) begin
      GEN_10 <= T_406_3_T_446_addr;
    end
    if(T_406_3_T_437_en & T_406_3_T_437_mask) begin
      T_406_3[T_406_3_T_437_addr] <= T_406_3_T_437_data;
    end
    if(T_406_4_T_446_en) begin
      GEN_13 <= T_406_4_T_446_addr;
    end
    if(T_406_4_T_437_en & T_406_4_T_437_mask) begin
      T_406_4[T_406_4_T_437_addr] <= T_406_4_T_437_data;
    end
    if(T_406_5_T_446_en) begin
      GEN_16 <= T_406_5_T_446_addr;
    end
    if(T_406_5_T_437_en & T_406_5_T_437_mask) begin
      T_406_5[T_406_5_T_437_addr] <= T_406_5_T_437_data;
    end
    if(T_406_6_T_446_en) begin
      GEN_19 <= T_406_6_T_446_addr;
    end
    if(T_406_6_T_437_en & T_406_6_T_437_mask) begin
      T_406_6[T_406_6_T_437_addr] <= T_406_6_T_437_data;
    end
    if(T_406_7_T_446_en) begin
      GEN_22 <= T_406_7_T_446_addr;
    end
    if(T_406_7_T_437_en & T_406_7_T_437_mask) begin
      T_406_7[T_406_7_T_437_addr] <= T_406_7_T_437_data;
    end
  end
endmodule
module Arbiter_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [11:0] io_in_0_bits_addr,
  input   io_in_0_bits_write,
  input  [63:0] io_in_0_bits_wdata,
  input  [7:0] io_in_0_bits_wmask,
  input   io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [11:0] io_in_1_bits_addr,
  input   io_in_1_bits_write,
  input  [63:0] io_in_1_bits_wdata,
  input  [7:0] io_in_1_bits_wmask,
  input   io_in_1_bits_way_en,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [11:0] io_in_2_bits_addr,
  input   io_in_2_bits_write,
  input  [63:0] io_in_2_bits_wdata,
  input  [7:0] io_in_2_bits_wmask,
  input   io_in_2_bits_way_en,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [11:0] io_in_3_bits_addr,
  input   io_in_3_bits_write,
  input  [63:0] io_in_3_bits_wdata,
  input  [7:0] io_in_3_bits_wmask,
  input   io_in_3_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [11:0] io_out_bits_addr,
  output  io_out_bits_write,
  output [63:0] io_out_bits_wdata,
  output [7:0] io_out_bits_wmask,
  output  io_out_bits_way_en,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [11:0] GEN_1;
  wire  GEN_2;
  wire [63:0] GEN_3;
  wire [7:0] GEN_4;
  wire  GEN_5;
  wire [1:0] GEN_6;
  wire [11:0] GEN_7;
  wire  GEN_8;
  wire [63:0] GEN_9;
  wire [7:0] GEN_10;
  wire  GEN_11;
  wire [1:0] GEN_12;
  wire [11:0] GEN_13;
  wire  GEN_14;
  wire [63:0] GEN_15;
  wire [7:0] GEN_16;
  wire  GEN_17;
  wire  T_2024;
  wire  T_2025;
  wire  grant_1;
  wire  grant_2;
  wire  grant_3;
  wire  T_2030;
  wire  T_2031;
  wire  T_2032;
  wire  T_2034;
  wire  T_2035;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_2030;
  assign io_in_2_ready = T_2031;
  assign io_in_3_ready = T_2032;
  assign io_out_valid = T_2035;
  assign io_out_bits_addr = GEN_13;
  assign io_out_bits_write = GEN_14;
  assign io_out_bits_wdata = GEN_15;
  assign io_out_bits_wmask = GEN_16;
  assign io_out_bits_way_en = GEN_17;
  assign io_chosen = GEN_12;
  assign GEN_0 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_1 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr;
  assign GEN_2 = io_in_2_valid ? io_in_2_bits_write : io_in_3_bits_write;
  assign GEN_3 = io_in_2_valid ? io_in_2_bits_wdata : io_in_3_bits_wdata;
  assign GEN_4 = io_in_2_valid ? io_in_2_bits_wmask : io_in_3_bits_wmask;
  assign GEN_5 = io_in_2_valid ? io_in_2_bits_way_en : io_in_3_bits_way_en;
  assign GEN_6 = io_in_1_valid ? 2'h1 : GEN_0;
  assign GEN_7 = io_in_1_valid ? io_in_1_bits_addr : GEN_1;
  assign GEN_8 = io_in_1_valid ? io_in_1_bits_write : GEN_2;
  assign GEN_9 = io_in_1_valid ? io_in_1_bits_wdata : GEN_3;
  assign GEN_10 = io_in_1_valid ? io_in_1_bits_wmask : GEN_4;
  assign GEN_11 = io_in_1_valid ? io_in_1_bits_way_en : GEN_5;
  assign GEN_12 = io_in_0_valid ? 2'h0 : GEN_6;
  assign GEN_13 = io_in_0_valid ? io_in_0_bits_addr : GEN_7;
  assign GEN_14 = io_in_0_valid ? io_in_0_bits_write : GEN_8;
  assign GEN_15 = io_in_0_valid ? io_in_0_bits_wdata : GEN_9;
  assign GEN_16 = io_in_0_valid ? io_in_0_bits_wmask : GEN_10;
  assign GEN_17 = io_in_0_valid ? io_in_0_bits_way_en : GEN_11;
  assign T_2024 = io_in_0_valid | io_in_1_valid;
  assign T_2025 = T_2024 | io_in_2_valid;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign grant_2 = T_2024 == 1'h0;
  assign grant_3 = T_2025 == 1'h0;
  assign T_2030 = grant_1 & io_out_ready;
  assign T_2031 = grant_2 & io_out_ready;
  assign T_2032 = grant_3 & io_out_ready;
  assign T_2034 = grant_3 == 1'h0;
  assign T_2035 = T_2034 | io_in_3_valid;
endmodule
module MetadataArray(
  input   clk,
  input   reset,
  output  io_read_ready,
  input   io_read_valid,
  input  [5:0] io_read_bits_idx,
  input   io_read_bits_way_en,
  output  io_write_ready,
  input   io_write_valid,
  input  [5:0] io_write_bits_idx,
  input   io_write_bits_way_en,
  input  [19:0] io_write_bits_data_tag,
  input  [1:0] io_write_bits_data_coh_state,
  output [19:0] io_resp_0_tag,
  output [1:0] io_resp_0_coh_state
);
  wire [1:0] T_44_state;
  wire [19:0] rstVal_tag;
  wire [1:0] rstVal_coh_state;
  reg [6:0] rst_cnt;
  reg [31:0] GEN_1;
  wire  rst;
  wire [6:0] waddr;
  wire [19:0] T_1569_tag;
  wire [1:0] T_1569_coh_state;
  wire [21:0] wdata;
  wire [7:0] T_1664;
  wire [6:0] T_1665;
  wire [6:0] GEN_0;
  reg [21:0] T_1674_0 [0:63];
  reg [31:0] GEN_2;
  wire [21:0] T_1674_0_T_1691_data;
  wire [5:0] T_1674_0_T_1691_addr;
  wire  T_1674_0_T_1691_en;
  reg [5:0] GEN_3;
  reg [31:0] GEN_4;
  wire [21:0] T_1674_0_T_1685_data;
  wire [5:0] T_1674_0_T_1685_addr;
  wire  T_1674_0_T_1685_mask;
  wire  T_1674_0_T_1685_en;
  wire  T_1675;
  wire [21:0] T_1681_0;
  wire [5:0] T_1688;
  wire [19:0] T_1777_tag;
  wire [1:0] T_1777_coh_state;
  wire [1:0] T_1861;
  wire [19:0] T_1862;
  wire  T_1864;
  wire  T_1866;
  wire  T_1867;
  assign io_read_ready = T_1867;
  assign io_write_ready = T_1864;
  assign io_resp_0_tag = T_1777_tag;
  assign io_resp_0_coh_state = T_1777_coh_state;
  assign T_44_state = 2'h0;
  assign rstVal_tag = 20'h0;
  assign rstVal_coh_state = T_44_state;
  assign rst = rst_cnt < 7'h40;
  assign waddr = rst ? rst_cnt : {{1'd0}, io_write_bits_idx};
  assign T_1569_tag = rst ? rstVal_tag : io_write_bits_data_tag;
  assign T_1569_coh_state = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign wdata = {T_1569_tag,T_1569_coh_state};
  assign T_1664 = rst_cnt + 7'h1;
  assign T_1665 = T_1664[6:0];
  assign GEN_0 = rst ? T_1665 : rst_cnt;
  assign T_1674_0_T_1691_addr = T_1688;
  assign T_1674_0_T_1691_en = io_read_valid;
  assign T_1674_0_T_1691_data = T_1674_0[GEN_3];
  assign T_1674_0_T_1685_data = T_1681_0;
  assign T_1674_0_T_1685_addr = waddr[5:0];
  assign T_1674_0_T_1685_mask = T_1675;
  assign T_1674_0_T_1685_en = T_1675;
  assign T_1675 = rst | io_write_valid;
  assign T_1681_0 = wdata;
  assign T_1688 = io_read_bits_idx;
  assign T_1777_tag = T_1862;
  assign T_1777_coh_state = T_1861;
  assign T_1861 = T_1674_0_T_1691_data[1:0];
  assign T_1862 = T_1674_0_T_1691_data[21:2];
  assign T_1864 = rst == 1'h0;
  assign T_1866 = io_write_valid == 1'h0;
  assign T_1867 = T_1864 & T_1866;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  rst_cnt = GEN_1[6:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_1674_0[initvar] = GEN_2[21:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {1{$random}};
  GEN_3 = GEN_4[5:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else begin
      if(rst) begin
        rst_cnt <= T_1665;
      end
    end
    if(T_1674_0_T_1691_en) begin
      GEN_3 <= T_1674_0_T_1691_addr;
    end
    if(T_1674_0_T_1685_en & T_1674_0_T_1685_mask) begin
      T_1674_0[T_1674_0_T_1685_addr] <= T_1674_0_T_1685_data;
    end
  end
endmodule
module AMOALU(
  input   clk,
  input   reset,
  input  [2:0] io_addr,
  input  [4:0] io_cmd,
  input  [1:0] io_typ,
  input  [63:0] io_lhs,
  input  [63:0] io_rhs,
  output [63:0] io_out
);
  wire  T_8;
  wire [31:0] T_9;
  wire [63:0] T_10;
  wire [63:0] rhs;
  wire  T_11;
  wire  T_12;
  wire  sgned;
  wire  T_14;
  wire  max;
  wire  T_16;
  wire  min;
  wire  T_19;
  wire [31:0] GEN_0;
  wire [31:0] T_20;
  wire [63:0] GEN_1;
  wire [63:0] T_21;
  wire [63:0] T_22;
  wire [63:0] T_23;
  wire [64:0] T_24;
  wire [63:0] adder_out;
  wire  T_25;
  wire  T_27;
  wire  T_30;
  wire  T_31;
  wire  T_32;
  wire  T_33;
  wire  T_34;
  wire  T_39;
  wire  T_40;
  wire  T_41;
  wire [31:0] T_42;
  wire [31:0] T_43;
  wire  T_44;
  wire [31:0] T_45;
  wire [31:0] T_46;
  wire  T_47;
  wire  T_50;
  wire  T_52;
  wire  T_53;
  wire  T_54;
  wire  T_55;
  wire  T_56;
  wire  T_57;
  wire  less;
  wire  T_58;
  wire  T_59;
  wire [63:0] T_60;
  wire  T_61;
  wire [63:0] T_62;
  wire  T_63;
  wire [63:0] T_64;
  wire  T_65;
  wire  T_67;
  wire [7:0] T_68;
  wire [15:0] T_69;
  wire [31:0] T_70;
  wire [63:0] T_71;
  wire  T_73;
  wire [15:0] T_74;
  wire [31:0] T_75;
  wire [63:0] T_76;
  wire [63:0] T_82;
  wire [63:0] T_83;
  wire [63:0] T_84;
  wire [63:0] T_85;
  wire [63:0] T_86;
  wire [63:0] T_87;
  wire [63:0] out;
  wire  T_89;
  wire  T_93;
  wire  T_97;
  wire  T_100;
  wire [1:0] T_101;
  wire  T_102;
  wire [1:0] T_104;
  wire  T_106;
  wire [1:0] T_109;
  wire [1:0] T_110;
  wire [1:0] T_113;
  wire [3:0] T_114;
  wire [3:0] T_117;
  wire  T_119;
  wire [3:0] T_122;
  wire [3:0] T_123;
  wire [3:0] T_126;
  wire [7:0] T_127;
  wire  T_128;
  wire  T_129;
  wire  T_130;
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire  T_134;
  wire  T_135;
  wire [7:0] T_139;
  wire [7:0] T_143;
  wire [7:0] T_147;
  wire [7:0] T_151;
  wire [7:0] T_155;
  wire [7:0] T_159;
  wire [7:0] T_163;
  wire [7:0] T_167;
  wire [15:0] T_168;
  wire [15:0] T_169;
  wire [31:0] T_170;
  wire [15:0] T_171;
  wire [15:0] T_172;
  wire [31:0] T_173;
  wire [63:0] wmask;
  wire [63:0] T_174;
  wire [63:0] T_175;
  wire [63:0] T_176;
  wire [63:0] T_177;
  assign io_out = T_177;
  assign T_8 = io_typ == 2'h2;
  assign T_9 = io_rhs[31:0];
  assign T_10 = {T_9,T_9};
  assign rhs = T_8 ? T_10 : io_rhs;
  assign T_11 = io_cmd == 5'hc;
  assign T_12 = io_cmd == 5'hd;
  assign sgned = T_11 | T_12;
  assign T_14 = io_cmd == 5'hf;
  assign max = T_12 | T_14;
  assign T_16 = io_cmd == 5'he;
  assign min = T_11 | T_16;
  assign T_19 = io_addr[2];
  assign GEN_0 = {{31'd0}, T_19};
  assign T_20 = GEN_0 << 31;
  assign GEN_1 = {{32'd0}, T_20};
  assign T_21 = 64'hffffffffffffffff ^ GEN_1;
  assign T_22 = io_lhs & T_21;
  assign T_23 = rhs & T_21;
  assign T_24 = T_22 + T_23;
  assign adder_out = T_24[63:0];
  assign T_25 = io_typ[0];
  assign T_27 = T_25 == 1'h0;
  assign T_30 = T_19 == 1'h0;
  assign T_31 = T_27 & T_30;
  assign T_32 = io_lhs[31];
  assign T_33 = io_lhs[63];
  assign T_34 = T_31 ? T_32 : T_33;
  assign T_39 = rhs[31];
  assign T_40 = rhs[63];
  assign T_41 = T_31 ? T_39 : T_40;
  assign T_42 = io_lhs[31:0];
  assign T_43 = rhs[31:0];
  assign T_44 = T_42 < T_43;
  assign T_45 = io_lhs[63:32];
  assign T_46 = rhs[63:32];
  assign T_47 = T_45 < T_46;
  assign T_50 = T_45 == T_46;
  assign T_52 = T_19 ? T_47 : T_44;
  assign T_53 = T_50 & T_44;
  assign T_54 = T_47 | T_53;
  assign T_55 = T_27 ? T_52 : T_54;
  assign T_56 = T_34 == T_41;
  assign T_57 = sgned ? T_34 : T_41;
  assign less = T_56 ? T_55 : T_57;
  assign T_58 = io_cmd == 5'h8;
  assign T_59 = io_cmd == 5'hb;
  assign T_60 = io_lhs & rhs;
  assign T_61 = io_cmd == 5'ha;
  assign T_62 = io_lhs | rhs;
  assign T_63 = io_cmd == 5'h9;
  assign T_64 = io_lhs ^ rhs;
  assign T_65 = less ? min : max;
  assign T_67 = io_typ == 2'h0;
  assign T_68 = io_rhs[7:0];
  assign T_69 = {T_68,T_68};
  assign T_70 = {T_69,T_69};
  assign T_71 = {T_70,T_70};
  assign T_73 = io_typ == 2'h1;
  assign T_74 = io_rhs[15:0];
  assign T_75 = {T_74,T_74};
  assign T_76 = {T_75,T_75};
  assign T_82 = T_73 ? T_76 : rhs;
  assign T_83 = T_67 ? T_71 : T_82;
  assign T_84 = T_65 ? io_lhs : T_83;
  assign T_85 = T_63 ? T_64 : T_84;
  assign T_86 = T_61 ? T_62 : T_85;
  assign T_87 = T_59 ? T_60 : T_86;
  assign out = T_58 ? adder_out : T_87;
  assign T_89 = io_addr[0];
  assign T_93 = io_typ >= 2'h1;
  assign T_97 = T_89 | T_93;
  assign T_100 = T_89 ? 1'h0 : 1'h1;
  assign T_101 = {T_97,T_100};
  assign T_102 = io_addr[1];
  assign T_104 = T_102 ? T_101 : 2'h0;
  assign T_106 = io_typ >= 2'h2;
  assign T_109 = T_106 ? 2'h3 : 2'h0;
  assign T_110 = T_104 | T_109;
  assign T_113 = T_102 ? 2'h0 : T_101;
  assign T_114 = {T_110,T_113};
  assign T_117 = T_19 ? T_114 : 4'h0;
  assign T_119 = io_typ >= 2'h3;
  assign T_122 = T_119 ? 4'hf : 4'h0;
  assign T_123 = T_117 | T_122;
  assign T_126 = T_19 ? 4'h0 : T_114;
  assign T_127 = {T_123,T_126};
  assign T_128 = T_127[0];
  assign T_129 = T_127[1];
  assign T_130 = T_127[2];
  assign T_131 = T_127[3];
  assign T_132 = T_127[4];
  assign T_133 = T_127[5];
  assign T_134 = T_127[6];
  assign T_135 = T_127[7];
  assign T_139 = T_128 ? 8'hff : 8'h0;
  assign T_143 = T_129 ? 8'hff : 8'h0;
  assign T_147 = T_130 ? 8'hff : 8'h0;
  assign T_151 = T_131 ? 8'hff : 8'h0;
  assign T_155 = T_132 ? 8'hff : 8'h0;
  assign T_159 = T_133 ? 8'hff : 8'h0;
  assign T_163 = T_134 ? 8'hff : 8'h0;
  assign T_167 = T_135 ? 8'hff : 8'h0;
  assign T_168 = {T_143,T_139};
  assign T_169 = {T_151,T_147};
  assign T_170 = {T_169,T_168};
  assign T_171 = {T_159,T_155};
  assign T_172 = {T_167,T_163};
  assign T_173 = {T_172,T_171};
  assign wmask = {T_173,T_170};
  assign T_174 = wmask & out;
  assign T_175 = ~ wmask;
  assign T_176 = T_175 & io_lhs;
  assign T_177 = T_174 | T_176;
endmodule
module DCache(
  input   clk,
  input   reset,
  output  io_cpu_req_ready,
  input   io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_addr,
  input  [5:0] io_cpu_req_bits_tag,
  input  [4:0] io_cpu_req_bits_cmd,
  input  [2:0] io_cpu_req_bits_typ,
  input   io_cpu_req_bits_phys,
  input  [63:0] io_cpu_req_bits_data,
  input   io_cpu_s1_kill,
  input  [63:0] io_cpu_s1_data,
  output  io_cpu_s2_nack,
  output  io_cpu_resp_valid,
  output [39:0] io_cpu_resp_bits_addr,
  output [5:0] io_cpu_resp_bits_tag,
  output [4:0] io_cpu_resp_bits_cmd,
  output [2:0] io_cpu_resp_bits_typ,
  output [63:0] io_cpu_resp_bits_data,
  output  io_cpu_resp_bits_replay,
  output  io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output [63:0] io_cpu_resp_bits_store_data,
  output  io_cpu_replay_next,
  output  io_cpu_xcpt_ma_ld,
  output  io_cpu_xcpt_ma_st,
  output  io_cpu_xcpt_pf_ld,
  output  io_cpu_xcpt_pf_st,
  input   io_cpu_invalidate_lr,
  output  io_cpu_ordered,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_pum,
  output  io_ptw_req_bits_mxr,
  output [26:0] io_ptw_req_bits_addr,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [15:0] io_ptw_resp_bits_pte_reserved_for_hardware,
  input  [37:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_a,
  input   io_ptw_resp_bits_pte_g,
  input   io_ptw_resp_bits_pte_u,
  input   io_ptw_resp_bits_pte_x,
  input   io_ptw_resp_bits_pte_w,
  input   io_ptw_resp_bits_pte_r,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [37:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [3:0] io_ptw_status_zero1,
  input   io_ptw_status_mxr,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output  io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [10:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_probe_ready,
  input   io_mem_probe_valid,
  input  [25:0] io_mem_probe_bits_addr_block,
  input  [1:0] io_mem_probe_bits_p_type,
  input   io_mem_release_ready,
  output  io_mem_release_valid,
  output [2:0] io_mem_release_bits_addr_beat,
  output [25:0] io_mem_release_bits_addr_block,
  output  io_mem_release_bits_client_xact_id,
  output  io_mem_release_bits_voluntary,
  output [2:0] io_mem_release_bits_r_type,
  output [63:0] io_mem_release_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input   io_mem_grant_bits_client_xact_id,
  input  [1:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [1:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id
);
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [1:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [1:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  wire  T_1924;
  reg [15:0] T_1927;
  reg [31:0] GEN_90;
  wire  T_1928;
  wire  T_1929;
  wire  T_1930;
  wire  T_1931;
  wire  T_1932;
  wire  T_1933;
  wire  T_1934;
  wire [14:0] T_1935;
  wire [15:0] T_1936;
  wire [15:0] GEN_2;
  wire  metaReadArb_clk;
  wire  metaReadArb_reset;
  wire  metaReadArb_io_in_0_ready;
  wire  metaReadArb_io_in_0_valid;
  wire [5:0] metaReadArb_io_in_0_bits_idx;
  wire  metaReadArb_io_in_0_bits_way_en;
  wire  metaReadArb_io_in_1_ready;
  wire  metaReadArb_io_in_1_valid;
  wire [5:0] metaReadArb_io_in_1_bits_idx;
  wire  metaReadArb_io_in_1_bits_way_en;
  wire  metaReadArb_io_in_2_ready;
  wire  metaReadArb_io_in_2_valid;
  wire [5:0] metaReadArb_io_in_2_bits_idx;
  wire  metaReadArb_io_in_2_bits_way_en;
  wire  metaReadArb_io_out_ready;
  wire  metaReadArb_io_out_valid;
  wire [5:0] metaReadArb_io_out_bits_idx;
  wire  metaReadArb_io_out_bits_way_en;
  wire [1:0] metaReadArb_io_chosen;
  wire  metaWriteArb_clk;
  wire  metaWriteArb_reset;
  wire  metaWriteArb_io_in_0_ready;
  wire  metaWriteArb_io_in_0_valid;
  wire [5:0] metaWriteArb_io_in_0_bits_idx;
  wire  metaWriteArb_io_in_0_bits_way_en;
  wire [19:0] metaWriteArb_io_in_0_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_0_bits_data_coh_state;
  wire  metaWriteArb_io_in_1_ready;
  wire  metaWriteArb_io_in_1_valid;
  wire [5:0] metaWriteArb_io_in_1_bits_idx;
  wire  metaWriteArb_io_in_1_bits_way_en;
  wire [19:0] metaWriteArb_io_in_1_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_1_bits_data_coh_state;
  wire  metaWriteArb_io_in_2_ready;
  wire  metaWriteArb_io_in_2_valid;
  wire [5:0] metaWriteArb_io_in_2_bits_idx;
  wire  metaWriteArb_io_in_2_bits_way_en;
  wire [19:0] metaWriteArb_io_in_2_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_2_bits_data_coh_state;
  wire  metaWriteArb_io_out_ready;
  wire  metaWriteArb_io_out_valid;
  wire [5:0] metaWriteArb_io_out_bits_idx;
  wire  metaWriteArb_io_out_bits_way_en;
  wire [19:0] metaWriteArb_io_out_bits_data_tag;
  wire [1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire [1:0] metaWriteArb_io_chosen;
  wire  data_clk;
  wire  data_reset;
  wire  data_io_req_valid;
  wire [11:0] data_io_req_bits_addr;
  wire  data_io_req_bits_write;
  wire [63:0] data_io_req_bits_wdata;
  wire [7:0] data_io_req_bits_wmask;
  wire  data_io_req_bits_way_en;
  wire [63:0] data_io_resp_0;
  wire  dataArb_clk;
  wire  dataArb_reset;
  wire  dataArb_io_in_0_ready;
  wire  dataArb_io_in_0_valid;
  wire [11:0] dataArb_io_in_0_bits_addr;
  wire  dataArb_io_in_0_bits_write;
  wire [63:0] dataArb_io_in_0_bits_wdata;
  wire [7:0] dataArb_io_in_0_bits_wmask;
  wire  dataArb_io_in_0_bits_way_en;
  wire  dataArb_io_in_1_ready;
  wire  dataArb_io_in_1_valid;
  wire [11:0] dataArb_io_in_1_bits_addr;
  wire  dataArb_io_in_1_bits_write;
  wire [63:0] dataArb_io_in_1_bits_wdata;
  wire [7:0] dataArb_io_in_1_bits_wmask;
  wire  dataArb_io_in_1_bits_way_en;
  wire  dataArb_io_in_2_ready;
  wire  dataArb_io_in_2_valid;
  wire [11:0] dataArb_io_in_2_bits_addr;
  wire  dataArb_io_in_2_bits_write;
  wire [63:0] dataArb_io_in_2_bits_wdata;
  wire [7:0] dataArb_io_in_2_bits_wmask;
  wire  dataArb_io_in_2_bits_way_en;
  wire  dataArb_io_in_3_ready;
  wire  dataArb_io_in_3_valid;
  wire [11:0] dataArb_io_in_3_bits_addr;
  wire  dataArb_io_in_3_bits_write;
  wire [63:0] dataArb_io_in_3_bits_wdata;
  wire [7:0] dataArb_io_in_3_bits_wmask;
  wire  dataArb_io_in_3_bits_way_en;
  wire  dataArb_io_out_ready;
  wire  dataArb_io_out_valid;
  wire [11:0] dataArb_io_out_bits_addr;
  wire  dataArb_io_out_bits_write;
  wire [63:0] dataArb_io_out_bits_wdata;
  wire [7:0] dataArb_io_out_bits_wmask;
  wire  dataArb_io_out_bits_way_en;
  wire [1:0] dataArb_io_chosen;
  wire  T_2218;
  reg  s1_valid;
  reg [31:0] GEN_91;
  wire  T_2220;
  reg  s1_probe;
  reg [31:0] GEN_95;
  reg [25:0] probe_bits_addr_block;
  reg [31:0] GEN_99;
  reg [1:0] probe_bits_p_type;
  reg [31:0] GEN_100;
  wire [25:0] GEN_3;
  wire [1:0] GEN_4;
  wire  s1_nack;
  wire  T_2247;
  wire  T_2248;
  wire [1:0] T_2249;
  wire [1:0] T_2250;
  wire [3:0] T_2251;
  wire  T_2253;
  wire  T_2255;
  wire  s1_valid_masked;
  wire  T_2257;
  wire  s1_valid_not_nacked;
  reg [39:0] s1_req_addr;
  reg [63:0] GEN_104;
  reg [5:0] s1_req_tag;
  reg [31:0] GEN_112;
  reg [4:0] s1_req_cmd;
  reg [31:0] GEN_121;
  reg [2:0] s1_req_typ;
  reg [31:0] GEN_132;
  reg  s1_req_phys;
  reg [31:0] GEN_133;
  reg [63:0] s1_req_data;
  reg [63:0] GEN_134;
  wire [27:0] T_2324;
  wire [5:0] T_2325;
  wire [33:0] T_2326;
  wire [39:0] T_2327;
  wire [39:0] GEN_5;
  wire [5:0] GEN_6;
  wire [4:0] GEN_7;
  wire [2:0] GEN_8;
  wire  GEN_9;
  wire [63:0] GEN_10;
  wire  T_2328;
  wire  T_2329;
  wire  T_2330;
  wire  T_2331;
  wire  T_2332;
  wire  T_2333;
  wire  T_2334;
  wire  T_2335;
  wire  s1_read;
  wire  T_2336;
  wire  T_2338;
  wire  s1_write;
  wire  s1_readwrite;
  reg  s1_flush_valid;
  reg [31:0] GEN_135;
  reg  grant_wait;
  reg [31:0] GEN_136;
  reg  release_ack_wait;
  reg [31:0] GEN_137;
  reg [2:0] release_state;
  reg [31:0] GEN_138;
  wire  pstore1_valid;
  reg  pstore2_valid;
  reg [31:0] GEN_139;
  wire  T_2348;
  wire  T_2349;
  wire  inWriteback;
  wire [1:0] releaseWay;
  wire  T_2351;
  wire  T_2353;
  wire  T_2354;
  wire  T_2357;
  wire  T_2358;
  wire  T_2359;
  wire  T_2360;
  wire  T_2361;
  wire  T_2362;
  wire  T_2363;
  wire  T_2364;
  wire  T_2365;
  wire  T_2366;
  wire  T_2367;
  wire  T_2372;
  wire  T_2382;
  wire  GEN_11;
  wire [5:0] T_2384;
  wire  T_2388;
  wire  GEN_12;
  wire  tlb_clk;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [27:0] tlb_io_req_bits_vpn;
  wire  tlb_io_req_bits_passthrough;
  wire  tlb_io_req_bits_instruction;
  wire  tlb_io_req_bits_store;
  wire  tlb_io_resp_miss;
  wire [19:0] tlb_io_resp_ppn;
  wire  tlb_io_resp_xcpt_ld;
  wire  tlb_io_resp_xcpt_st;
  wire  tlb_io_resp_xcpt_if;
  wire  tlb_io_resp_cacheable;
  wire  tlb_io_ptw_req_ready;
  wire  tlb_io_ptw_req_valid;
  wire [1:0] tlb_io_ptw_req_bits_prv;
  wire  tlb_io_ptw_req_bits_pum;
  wire  tlb_io_ptw_req_bits_mxr;
  wire [26:0] tlb_io_ptw_req_bits_addr;
  wire  tlb_io_ptw_req_bits_store;
  wire  tlb_io_ptw_req_bits_fetch;
  wire  tlb_io_ptw_resp_valid;
  wire [15:0] tlb_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] tlb_io_ptw_resp_bits_pte_ppn;
  wire [1:0] tlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  tlb_io_ptw_resp_bits_pte_d;
  wire  tlb_io_ptw_resp_bits_pte_a;
  wire  tlb_io_ptw_resp_bits_pte_g;
  wire  tlb_io_ptw_resp_bits_pte_u;
  wire  tlb_io_ptw_resp_bits_pte_x;
  wire  tlb_io_ptw_resp_bits_pte_w;
  wire  tlb_io_ptw_resp_bits_pte_r;
  wire  tlb_io_ptw_resp_bits_pte_v;
  wire [6:0] tlb_io_ptw_ptbr_asid;
  wire [37:0] tlb_io_ptw_ptbr_ppn;
  wire  tlb_io_ptw_invalidate;
  wire  tlb_io_ptw_status_debug;
  wire [1:0] tlb_io_ptw_status_prv;
  wire  tlb_io_ptw_status_sd;
  wire [30:0] tlb_io_ptw_status_zero3;
  wire  tlb_io_ptw_status_sd_rv32;
  wire [1:0] tlb_io_ptw_status_zero2;
  wire [4:0] tlb_io_ptw_status_vm;
  wire [3:0] tlb_io_ptw_status_zero1;
  wire  tlb_io_ptw_status_mxr;
  wire  tlb_io_ptw_status_pum;
  wire  tlb_io_ptw_status_mprv;
  wire [1:0] tlb_io_ptw_status_xs;
  wire [1:0] tlb_io_ptw_status_fs;
  wire [1:0] tlb_io_ptw_status_mpp;
  wire [1:0] tlb_io_ptw_status_hpp;
  wire  tlb_io_ptw_status_spp;
  wire  tlb_io_ptw_status_mpie;
  wire  tlb_io_ptw_status_hpie;
  wire  tlb_io_ptw_status_spie;
  wire  tlb_io_ptw_status_upie;
  wire  tlb_io_ptw_status_mie;
  wire  tlb_io_ptw_status_hie;
  wire  tlb_io_ptw_status_sie;
  wire  tlb_io_ptw_status_uie;
  wire  T_2390;
  wire [27:0] T_2391;
  wire  T_2394;
  wire  T_2396;
  wire  T_2397;
  wire  GEN_13;
  wire  T_2399;
  wire  T_2400;
  wire [11:0] T_2402;
  wire [31:0] s1_paddr;
  wire [19:0] T_2403;
  wire [19:0] T_2404;
  wire [19:0] s1_tag;
  wire  s1_victim_way;
  wire  MetadataArray_1_clk;
  wire  MetadataArray_1_reset;
  wire  MetadataArray_1_io_read_ready;
  wire  MetadataArray_1_io_read_valid;
  wire [5:0] MetadataArray_1_io_read_bits_idx;
  wire  MetadataArray_1_io_read_bits_way_en;
  wire  MetadataArray_1_io_write_ready;
  wire  MetadataArray_1_io_write_valid;
  wire [5:0] MetadataArray_1_io_write_bits_idx;
  wire  MetadataArray_1_io_write_bits_way_en;
  wire [19:0] MetadataArray_1_io_write_bits_data_tag;
  wire [1:0] MetadataArray_1_io_write_bits_data_coh_state;
  wire [19:0] MetadataArray_1_io_resp_0_tag;
  wire [1:0] MetadataArray_1_io_resp_0_coh_state;
  wire  T_2406;
  wire  T_2407;
  wire  s1_hit_way;
  wire [1:0] T_2431_state;
  wire [1:0] T_2455;
  wire [1:0] s1_hit_state_state;
  reg  s2_valid;
  reg [31:0] GEN_140;
  reg  s2_probe;
  reg [31:0] GEN_141;
  wire  T_2587;
  wire  T_2588;
  wire  releaseInFlight;
  reg  T_2591;
  reg [31:0] GEN_142;
  wire  s2_valid_masked;
  reg [39:0] s2_req_addr;
  reg [63:0] GEN_143;
  reg [5:0] s2_req_tag;
  reg [31:0] GEN_144;
  reg [4:0] s2_req_cmd;
  reg [31:0] GEN_145;
  reg [2:0] s2_req_typ;
  reg [31:0] GEN_146;
  reg  s2_req_phys;
  reg [31:0] GEN_147;
  reg [63:0] s2_req_data;
  reg [63:0] GEN_148;
  reg  s2_uncached;
  reg [31:0] GEN_149;
  wire  T_2659;
  wire  T_2661;
  wire [39:0] GEN_15;
  wire [5:0] GEN_16;
  wire [4:0] GEN_17;
  wire [2:0] GEN_18;
  wire  GEN_19;
  wire [63:0] GEN_20;
  wire  GEN_21;
  wire  T_2664;
  wire  T_2665;
  wire  T_2666;
  wire  T_2667;
  wire  T_2668;
  wire  T_2669;
  wire  T_2670;
  wire  T_2671;
  wire  s2_read;
  wire  T_2672;
  wire  T_2674;
  wire  s2_write;
  wire  s2_readwrite;
  reg  s2_flush_valid;
  reg [31:0] GEN_150;
  wire  T_2678;
  reg [63:0] s2_data;
  reg [63:0] GEN_151;
  wire [63:0] GEN_22;
  reg  s2_probe_way;
  reg [31:0] GEN_152;
  wire  GEN_23;
  reg [1:0] s2_probe_state_state;
  reg [31:0] GEN_153;
  wire [1:0] GEN_24;
  reg  s2_hit_way;
  reg [31:0] GEN_154;
  wire  GEN_25;
  reg [1:0] s2_hit_state_state;
  reg [31:0] GEN_155;
  wire [1:0] GEN_26;
  wire  T_2728;
  wire  T_2729;
  wire  T_2731;
  wire  T_2732;
  wire  T_2733;
  wire  T_2734;
  wire  s2_hit;
  wire  T_2738;
  wire  s2_valid_hit;
  wire  T_2741;
  wire  T_2742;
  wire  T_2743;
  wire  T_2745;
  wire  T_2746;
  wire  T_2748;
  wire  s2_valid_miss;
  wire  T_2750;
  wire  s2_valid_cached_miss;
  wire  s2_victimize;
  wire  s2_valid_uncached;
  wire  T_2751;
  wire  T_2753;
  wire  T_2754;
  reg  T_2756;
  reg [31:0] GEN_156;
  wire  GEN_27;
  wire [1:0] T_2758;
  wire [1:0] s2_victim_way;
  reg [19:0] s2_victim_tag;
  reg [31:0] GEN_157;
  wire [19:0] GEN_0_tag;
  wire [1:0] GEN_0_coh_state;
  wire [19:0] GEN_28;
  wire [1:0] GEN_29;
  wire [19:0] GEN_30;
  reg [1:0] T_2766_state;
  reg [31:0] GEN_158;
  wire [19:0] GEN_1_tag;
  wire [1:0] GEN_1_coh_state;
  wire [1:0] GEN_33;
  wire [1:0] s2_victim_state_state;
  wire  s2_victim_dirty;
  wire [1:0] T_2816;
  wire [1:0] s2_new_hit_state_state;
  wire  T_2860;
  wire  s2_update_meta;
  wire  T_2863;
  wire  T_2864;
  wire  T_2865;
  wire  T_2867;
  wire  T_2868;
  wire  T_2871;
  wire  T_2872;
  wire  GEN_34;
  wire [1:0] T_2875;
  wire [3:0] T_2877;
  wire [4:0] T_2879;
  wire [3:0] T_2880;
  wire [2:0] T_2881;
  wire [39:0] GEN_0;
  wire [39:0] T_2882;
  wire  misaligned;
  wire  T_2884;
  wire  T_2885;
  wire  T_2886;
  wire  T_2887;
  reg [4:0] lrscCount;
  reg [31:0] GEN_159;
  wire  lrscValid;
  reg [33:0] lrscAddr;
  reg [63:0] GEN_160;
  wire [33:0] T_2895;
  wire  T_2896;
  wire  T_2897;
  wire  T_2899;
  wire  s2_sc_fail;
  wire  T_2900;
  wire [4:0] GEN_35;
  wire [33:0] GEN_36;
  wire [5:0] T_2904;
  wire [4:0] T_2905;
  wire [4:0] GEN_37;
  wire  T_2906;
  wire  T_2907;
  wire [4:0] GEN_38;
  wire  T_2909;
  reg [4:0] pstore1_cmd;
  reg [31:0] GEN_161;
  wire [4:0] GEN_39;
  reg [2:0] pstore1_typ;
  reg [31:0] GEN_162;
  wire [2:0] GEN_40;
  reg [31:0] pstore1_addr;
  reg [31:0] GEN_163;
  wire [31:0] GEN_41;
  reg [63:0] pstore1_data;
  reg [63:0] GEN_164;
  wire [63:0] GEN_42;
  reg  pstore1_way;
  reg [31:0] GEN_165;
  wire  GEN_43;
  wire [1:0] T_2914;
  wire  T_2916;
  wire [7:0] T_2917;
  wire [15:0] T_2918;
  wire [31:0] T_2919;
  wire [63:0] T_2920;
  wire  T_2922;
  wire [15:0] T_2923;
  wire [31:0] T_2924;
  wire [63:0] T_2925;
  wire  T_2927;
  wire [31:0] T_2928;
  wire [63:0] T_2929;
  wire [63:0] T_2930;
  wire [63:0] T_2931;
  wire [63:0] T_2932;
  wire [63:0] pstore1_storegen_data;
  wire  T_2934;
  wire  T_2935;
  wire  T_2936;
  wire  T_2937;
  wire  T_2938;
  wire  T_2939;
  wire  T_2940;
  wire  T_2941;
  wire  T_2942;
  wire  T_2943;
  wire  T_2944;
  wire  T_2945;
  wire  pstore_drain_structural;
  wire  pstore_drain_opportunistic;
  wire  pstore_drain_on_miss;
  wire  T_2960;
  wire  T_2961;
  wire  T_2962;
  wire  T_2963;
  wire  T_2964;
  wire  pstore_drain;
  wire  T_2965;
  wire  T_2967;
  wire  T_2968;
  reg  T_2970;
  reg [31:0] GEN_166;
  wire  T_2972;
  wire  T_2974;
  wire  T_2975;
  wire  T_2976;
  wire  T_2978;
  wire  T_2979;
  wire  T_2980;
  wire  T_2982;
  wire  T_2983;
  wire  T_2985;
  wire  advance_pstore1;
  wire  T_2988;
  wire  T_2989;
  reg [31:0] pstore2_addr;
  reg [31:0] GEN_167;
  wire [31:0] GEN_44;
  reg  pstore2_way;
  reg [31:0] GEN_168;
  wire  GEN_45;
  reg [63:0] pstore2_storegen_data;
  reg [63:0] GEN_169;
  wire [63:0] GEN_46;
  wire  T_2991;
  wire  T_2995;
  wire  T_2999;
  wire  T_3002;
  wire [1:0] T_3003;
  wire  T_3004;
  wire [1:0] T_3006;
  wire  T_3008;
  wire [1:0] T_3011;
  wire [1:0] T_3012;
  wire [1:0] T_3015;
  wire [3:0] T_3016;
  wire  T_3017;
  wire [3:0] T_3019;
  wire  T_3021;
  wire [3:0] T_3024;
  wire [3:0] T_3025;
  wire [3:0] T_3028;
  wire [7:0] T_3029;
  reg [7:0] pstore2_storegen_mask;
  reg [31:0] GEN_170;
  wire [7:0] GEN_47;
  wire [31:0] T_3031;
  wire  T_3032;
  wire [63:0] T_3033;
  wire [7:0] T_3076;
  wire [22:0] GEN_1;
  wire [22:0] T_3077;
  wire [8:0] s1_idx;
  wire [8:0] T_3078;
  wire  T_3079;
  wire  T_3080;
  wire [8:0] T_3081;
  wire  T_3082;
  wire  T_3083;
  wire  T_3084;
  wire  s1_raw_hazard;
  wire  T_3085;
  wire  GEN_48;
  wire  T_3087;
  wire  T_3089;
  wire  T_3090;
  wire  T_3091;
  wire [5:0] T_3092;
  wire [1:0] T_3116_state;
  wire [1:0] T_3138_state;
  wire [19:0] T_3160;
  wire [25:0] T_3162;
  wire [5:0] T_3177;
  wire [25:0] cachedGetMessage_addr_block;
  wire  cachedGetMessage_client_xact_id;
  wire [2:0] cachedGetMessage_addr_beat;
  wire  cachedGetMessage_is_builtin_type;
  wire [2:0] cachedGetMessage_a_type;
  wire [10:0] cachedGetMessage_union;
  wire [63:0] cachedGetMessage_data;
  wire [2:0] T_3237;
  wire [2:0] T_3238;
  wire [1:0] T_3269;
  wire [4:0] T_3279;
  wire [10:0] T_3280;
  wire [25:0] uncachedGetMessage_addr_block;
  wire  uncachedGetMessage_client_xact_id;
  wire [2:0] uncachedGetMessage_addr_beat;
  wire  uncachedGetMessage_is_builtin_type;
  wire [2:0] uncachedGetMessage_a_type;
  wire [10:0] uncachedGetMessage_union;
  wire [63:0] uncachedGetMessage_data;
  wire [22:0] GEN_125;
  wire [22:0] T_3427;
  wire [7:0] T_3465;
  wire [8:0] T_3475;
  wire [10:0] T_3495;
  wire [25:0] uncachedPutMessage_addr_block;
  wire  uncachedPutMessage_client_xact_id;
  wire [2:0] uncachedPutMessage_addr_beat;
  wire  uncachedPutMessage_is_builtin_type;
  wire [2:0] uncachedPutMessage_a_type;
  wire [10:0] uncachedPutMessage_union;
  wire [63:0] uncachedPutMessage_data;
  wire [10:0] T_3617;
  wire [25:0] uncachedPutAtomicMessage_addr_block;
  wire  uncachedPutAtomicMessage_client_xact_id;
  wire [2:0] uncachedPutAtomicMessage_addr_beat;
  wire  uncachedPutAtomicMessage_is_builtin_type;
  wire [2:0] uncachedPutAtomicMessage_a_type;
  wire [10:0] uncachedPutAtomicMessage_union;
  wire [63:0] uncachedPutAtomicMessage_data;
  wire  T_3704;
  wire  T_3705;
  wire  T_3706;
  wire  T_3708;
  wire  T_3711;
  wire  T_3712;
  wire  T_3713;
  wire  T_3715;
  wire [25:0] GEN_49;
  wire  GEN_50;
  wire [2:0] GEN_51;
  wire  GEN_52;
  wire [2:0] GEN_53;
  wire [10:0] GEN_54;
  wire [63:0] GEN_55;
  wire [25:0] GEN_56;
  wire  GEN_57;
  wire [2:0] GEN_58;
  wire  GEN_59;
  wire [2:0] GEN_60;
  wire [10:0] GEN_61;
  wire [63:0] GEN_62;
  wire [25:0] GEN_63;
  wire  GEN_64;
  wire [2:0] GEN_65;
  wire  GEN_66;
  wire [2:0] GEN_67;
  wire [10:0] GEN_68;
  wire [63:0] GEN_69;
  wire  T_3716;
  wire  GEN_70;
  wire [2:0] T_3725_0;
  wire [3:0] GEN_126;
  wire  T_3727;
  wire  T_3728;
  wire  T_3729;
  wire  grantIsVoluntary;
  wire  T_3733;
  wire  T_3735;
  wire  grantIsUncached;
  wire  T_3736;
  wire  T_3737;
  wire  T_3738;
  wire  T_3740;
  wire [63:0] GEN_71;
  wire  GEN_72;
  wire [63:0] GEN_73;
  wire  GEN_74;
  wire  T_3742;
  wire  T_3743;
  reg [2:0] refillCount;
  reg [31:0] GEN_171;
  wire  T_3746;
  wire [3:0] T_3748;
  wire [2:0] T_3749;
  wire [2:0] GEN_75;
  wire  refillDone;
  wire  grantDone;
  wire  T_3751;
  wire  GEN_76;
  wire  T_3753;
  wire  T_3756;
  wire  T_3757;
  wire  T_3758;
  wire  T_3760;
  wire [28:0] T_3763;
  wire [31:0] GEN_127;
  wire [31:0] T_3764;
  wire  T_3768;
  wire  T_3769;
  wire  T_3770;
  wire  T_3772;
  wire [1:0] T_3781;
  wire [1:0] T_3782;
  wire [1:0] T_3805_state;
  wire  T_3838;
  wire  T_3841;
  wire  T_3842;
  wire [1:0] T_3866_manager_xact_id;
  wire  T_3866_manager_id;
  wire  T_3889;
  wire  T_3891;
  wire  T_3893;
  wire  block_probe;
  wire  T_3896;
  wire  T_3897;
  wire  T_3900;
  wire  T_3902;
  wire  T_3903;
  wire  T_3905;
  wire  T_3906;
  wire  T_3907;
  wire  T_3910;
  wire  T_3911;
  reg [2:0] writebackCount;
  reg [31:0] GEN_172;
  wire  T_3914;
  wire [3:0] T_3916;
  wire [2:0] T_3917;
  wire [2:0] GEN_78;
  wire  writebackDone;
  wire  T_3920;
  wire  T_3921;
  wire  releaseDone;
  wire  T_3923;
  wire  releaseRejected;
  wire  T_3924;
  reg  s1_release_data_valid;
  reg [31:0] GEN_173;
  wire  T_3926;
  wire  T_3927;
  reg  s2_release_data_valid;
  reg [31:0] GEN_174;
  wire [3:0] T_3929;
  wire [1:0] T_3932;
  wire [1:0] GEN_128;
  wire [2:0] T_3933;
  wire [1:0] T_3934;
  wire [1:0] T_3935;
  wire [3:0] GEN_129;
  wire [4:0] T_3936;
  wire [3:0] releaseDataBeat;
  wire [1:0] T_3960_state;
  wire  T_3985;
  wire [2:0] T_3986;
  wire  T_4015;
  wire [2:0] T_4016;
  wire  T_4017;
  wire [2:0] T_4018;
  wire  T_4019;
  wire [2:0] T_4020;
  wire [2:0] T_4049_addr_beat;
  wire [25:0] T_4049_addr_block;
  wire  T_4049_client_xact_id;
  wire  T_4049_voluntary;
  wire [2:0] T_4049_r_type;
  wire [63:0] T_4049_data;
  wire [2:0] T_4082;
  wire [2:0] voluntaryReleaseMessage_addr_beat;
  wire [25:0] voluntaryReleaseMessage_addr_block;
  wire  voluntaryReleaseMessage_client_xact_id;
  wire  voluntaryReleaseMessage_voluntary;
  wire [2:0] voluntaryReleaseMessage_r_type;
  wire [63:0] voluntaryReleaseMessage_data;
  wire [1:0] voluntaryNewCoh_state;
  wire  T_4196;
  wire [2:0] T_4197;
  wire [2:0] T_4227;
  wire [2:0] T_4229;
  wire [2:0] T_4231;
  wire [2:0] probeResponseMessage_addr_beat;
  wire [25:0] probeResponseMessage_addr_block;
  wire  probeResponseMessage_client_xact_id;
  wire  probeResponseMessage_voluntary;
  wire [2:0] probeResponseMessage_r_type;
  wire [63:0] probeResponseMessage_data;
  wire [1:0] T_4287;
  wire [1:0] T_4289;
  wire [1:0] T_4291;
  wire [1:0] probeNewCoh_state;
  wire [1:0] newCoh_state;
  wire  T_4356;
  wire  T_4358;
  wire  T_4360;
  wire  T_4361;
  wire  T_4363;
  wire [25:0] T_4365;
  wire [2:0] GEN_79;
  wire [25:0] GEN_80;
  wire [2:0] GEN_81;
  wire  T_4367;
  wire  T_4369;
  wire  T_4370;
  wire [2:0] GEN_82;
  wire  T_4374;
  wire  T_4375;
  wire  GEN_83;
  wire [2:0] GEN_84;
  wire [2:0] GEN_85;
  wire  GEN_86;
  wire [2:0] GEN_87;
  wire  T_4377;
  wire  T_4378;
  wire  T_4379;
  wire  GEN_88;
  wire  T_4383;
  wire [2:0] GEN_89;
  wire  GEN_92;
  wire  GEN_93;
  wire [2:0] GEN_94;
  wire [2:0] GEN_96;
  wire  T_4385;
  wire  T_4386;
  wire [2:0] GEN_97;
  wire  GEN_98;
  wire  GEN_101;
  wire  GEN_102;
  wire [2:0] GEN_103;
  wire [1:0] GEN_105;
  wire [1:0] GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire  T_4390;
  wire  T_4391;
  wire  GEN_109;
  wire  T_4394;
  wire  T_4395;
  wire [2:0] T_4397;
  wire [28:0] T_4398;
  wire [31:0] GEN_130;
  wire [31:0] T_4399;
  wire  T_4403;
  wire  T_4404;
  wire [28:0] T_4406;
  wire [31:0] T_4407;
  wire [5:0] T_4408;
  wire [19:0] T_4412;
  wire  T_4413;
  wire [2:0] GEN_110;
  wire  T_4415;
  wire  T_4416;
  wire  T_4418;
  wire  T_4419;
  reg  doUncachedResp;
  reg [31:0] GEN_175;
  wire  T_4422;
  wire  T_4424;
  wire  GEN_111;
  wire [63:0] s2_data_word;
  wire  T_4429;
  wire  T_4431;
  wire  T_4433;
  wire [31:0] T_4434;
  wire [31:0] T_4435;
  wire [31:0] T_4436;
  wire  T_4442;
  wire  T_4444;
  wire  T_4445;
  wire [31:0] T_4449;
  wire [31:0] T_4451;
  wire [63:0] T_4452;
  wire  T_4453;
  wire [15:0] T_4454;
  wire [15:0] T_4455;
  wire [15:0] T_4456;
  wire  T_4462;
  wire  T_4464;
  wire  T_4465;
  wire [47:0] T_4469;
  wire [47:0] T_4470;
  wire [47:0] T_4471;
  wire [63:0] T_4472;
  wire  T_4473;
  wire [7:0] T_4474;
  wire [7:0] T_4475;
  wire [7:0] T_4476;
  wire [7:0] T_4480;
  wire  T_4482;
  wire  T_4483;
  wire  T_4484;
  wire  T_4485;
  wire [55:0] T_4489;
  wire [55:0] T_4490;
  wire [55:0] T_4491;
  wire [63:0] T_4492;
  wire [63:0] GEN_131;
  wire [63:0] T_4493;
  wire  AMOALU_1_clk;
  wire  AMOALU_1_reset;
  wire [2:0] AMOALU_1_io_addr;
  wire [4:0] AMOALU_1_io_cmd;
  wire [1:0] AMOALU_1_io_typ;
  wire [63:0] AMOALU_1_io_lhs;
  wire [63:0] AMOALU_1_io_rhs;
  wire [63:0] AMOALU_1_io_out;
  reg  flushed;
  reg [31:0] GEN_176;
  reg  flushing;
  reg [31:0] GEN_177;
  reg [5:0] T_4517;
  reg [31:0] GEN_178;
  wire  T_4521;
  wire  GEN_113;
  wire  T_4523;
  wire  T_4524;
  wire  T_4526;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  T_4531;
  wire  T_4533;
  wire  T_4534;
  wire  T_4537;
  wire  T_4539;
  wire  T_4542;
  wire  T_4547;
  wire [6:0] T_4549;
  wire [5:0] T_4550;
  wire  GEN_117;
  wire [5:0] GEN_118;
  wire  GEN_119;
  wire  T_4553;
  wire  T_4556;
  wire  GEN_120;
  wire [5:0] GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire [63:0] GEN_14;
  reg [63:0] GEN_179;
  wire [7:0] GEN_31;
  reg [31:0] GEN_180;
  wire [63:0] GEN_32;
  reg [63:0] GEN_181;
  wire [7:0] GEN_77;
  reg [31:0] GEN_182;
  FinishQueue fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  Arbiter metaReadArb (
    .clk(metaReadArb_clk),
    .reset(metaReadArb_reset),
    .io_in_0_ready(metaReadArb_io_in_0_ready),
    .io_in_0_valid(metaReadArb_io_in_0_valid),
    .io_in_0_bits_idx(metaReadArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaReadArb_io_in_0_bits_way_en),
    .io_in_1_ready(metaReadArb_io_in_1_ready),
    .io_in_1_valid(metaReadArb_io_in_1_valid),
    .io_in_1_bits_idx(metaReadArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaReadArb_io_in_1_bits_way_en),
    .io_in_2_ready(metaReadArb_io_in_2_ready),
    .io_in_2_valid(metaReadArb_io_in_2_valid),
    .io_in_2_bits_idx(metaReadArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaReadArb_io_in_2_bits_way_en),
    .io_out_ready(metaReadArb_io_out_ready),
    .io_out_valid(metaReadArb_io_out_valid),
    .io_out_bits_idx(metaReadArb_io_out_bits_idx),
    .io_out_bits_way_en(metaReadArb_io_out_bits_way_en),
    .io_chosen(metaReadArb_io_chosen)
  );
  Arbiter_1 metaWriteArb (
    .clk(metaWriteArb_clk),
    .reset(metaWriteArb_reset),
    .io_in_0_ready(metaWriteArb_io_in_0_ready),
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_idx(metaWriteArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaWriteArb_io_in_0_bits_way_en),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_coh_state(metaWriteArb_io_in_0_bits_data_coh_state),
    .io_in_1_ready(metaWriteArb_io_in_1_ready),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_idx(metaWriteArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaWriteArb_io_in_1_bits_way_en),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_coh_state(metaWriteArb_io_in_1_bits_data_coh_state),
    .io_in_2_ready(metaWriteArb_io_in_2_ready),
    .io_in_2_valid(metaWriteArb_io_in_2_valid),
    .io_in_2_bits_idx(metaWriteArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaWriteArb_io_in_2_bits_way_en),
    .io_in_2_bits_data_tag(metaWriteArb_io_in_2_bits_data_tag),
    .io_in_2_bits_data_coh_state(metaWriteArb_io_in_2_bits_data_coh_state),
    .io_out_ready(metaWriteArb_io_out_ready),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_idx(metaWriteArb_io_out_bits_idx),
    .io_out_bits_way_en(metaWriteArb_io_out_bits_way_en),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_coh_state(metaWriteArb_io_out_bits_data_coh_state),
    .io_chosen(metaWriteArb_io_chosen)
  );
  DCacheDataArray data (
    .clk(data_clk),
    .reset(data_reset),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_wmask(data_io_req_bits_wmask),
    .io_req_bits_way_en(data_io_req_bits_way_en),
    .io_resp_0(data_io_resp_0)
  );
  Arbiter_2 dataArb (
    .clk(dataArb_clk),
    .reset(dataArb_reset),
    .io_in_0_ready(dataArb_io_in_0_ready),
    .io_in_0_valid(dataArb_io_in_0_valid),
    .io_in_0_bits_addr(dataArb_io_in_0_bits_addr),
    .io_in_0_bits_write(dataArb_io_in_0_bits_write),
    .io_in_0_bits_wdata(dataArb_io_in_0_bits_wdata),
    .io_in_0_bits_wmask(dataArb_io_in_0_bits_wmask),
    .io_in_0_bits_way_en(dataArb_io_in_0_bits_way_en),
    .io_in_1_ready(dataArb_io_in_1_ready),
    .io_in_1_valid(dataArb_io_in_1_valid),
    .io_in_1_bits_addr(dataArb_io_in_1_bits_addr),
    .io_in_1_bits_write(dataArb_io_in_1_bits_write),
    .io_in_1_bits_wdata(dataArb_io_in_1_bits_wdata),
    .io_in_1_bits_wmask(dataArb_io_in_1_bits_wmask),
    .io_in_1_bits_way_en(dataArb_io_in_1_bits_way_en),
    .io_in_2_ready(dataArb_io_in_2_ready),
    .io_in_2_valid(dataArb_io_in_2_valid),
    .io_in_2_bits_addr(dataArb_io_in_2_bits_addr),
    .io_in_2_bits_write(dataArb_io_in_2_bits_write),
    .io_in_2_bits_wdata(dataArb_io_in_2_bits_wdata),
    .io_in_2_bits_wmask(dataArb_io_in_2_bits_wmask),
    .io_in_2_bits_way_en(dataArb_io_in_2_bits_way_en),
    .io_in_3_ready(dataArb_io_in_3_ready),
    .io_in_3_valid(dataArb_io_in_3_valid),
    .io_in_3_bits_addr(dataArb_io_in_3_bits_addr),
    .io_in_3_bits_write(dataArb_io_in_3_bits_write),
    .io_in_3_bits_wdata(dataArb_io_in_3_bits_wdata),
    .io_in_3_bits_wmask(dataArb_io_in_3_bits_wmask),
    .io_in_3_bits_way_en(dataArb_io_in_3_bits_way_en),
    .io_out_ready(dataArb_io_out_ready),
    .io_out_valid(dataArb_io_out_valid),
    .io_out_bits_addr(dataArb_io_out_bits_addr),
    .io_out_bits_write(dataArb_io_out_bits_write),
    .io_out_bits_wdata(dataArb_io_out_bits_wdata),
    .io_out_bits_wmask(dataArb_io_out_bits_wmask),
    .io_out_bits_way_en(dataArb_io_out_bits_way_en),
    .io_chosen(dataArb_io_chosen)
  );
  TLB tlb (
    .clk(tlb_clk),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vpn(tlb_io_req_bits_vpn),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_instruction(tlb_io_req_bits_instruction),
    .io_req_bits_store(tlb_io_req_bits_store),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_ppn(tlb_io_resp_ppn),
    .io_resp_xcpt_ld(tlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(tlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(tlb_io_resp_xcpt_if),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_prv(tlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(tlb_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(tlb_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(tlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(tlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(tlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(tlb_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(tlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(tlb_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(tlb_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(tlb_io_ptw_invalidate),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_status_sd(tlb_io_ptw_status_sd),
    .io_ptw_status_zero3(tlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(tlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(tlb_io_ptw_status_zero2),
    .io_ptw_status_vm(tlb_io_ptw_status_vm),
    .io_ptw_status_zero1(tlb_io_ptw_status_zero1),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_pum(tlb_io_ptw_status_pum),
    .io_ptw_status_mprv(tlb_io_ptw_status_mprv),
    .io_ptw_status_xs(tlb_io_ptw_status_xs),
    .io_ptw_status_fs(tlb_io_ptw_status_fs),
    .io_ptw_status_mpp(tlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(tlb_io_ptw_status_hpp),
    .io_ptw_status_spp(tlb_io_ptw_status_spp),
    .io_ptw_status_mpie(tlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(tlb_io_ptw_status_hpie),
    .io_ptw_status_spie(tlb_io_ptw_status_spie),
    .io_ptw_status_upie(tlb_io_ptw_status_upie),
    .io_ptw_status_mie(tlb_io_ptw_status_mie),
    .io_ptw_status_hie(tlb_io_ptw_status_hie),
    .io_ptw_status_sie(tlb_io_ptw_status_sie),
    .io_ptw_status_uie(tlb_io_ptw_status_uie)
  );
  MetadataArray MetadataArray_1 (
    .clk(MetadataArray_1_clk),
    .reset(MetadataArray_1_reset),
    .io_read_ready(MetadataArray_1_io_read_ready),
    .io_read_valid(MetadataArray_1_io_read_valid),
    .io_read_bits_idx(MetadataArray_1_io_read_bits_idx),
    .io_read_bits_way_en(MetadataArray_1_io_read_bits_way_en),
    .io_write_ready(MetadataArray_1_io_write_ready),
    .io_write_valid(MetadataArray_1_io_write_valid),
    .io_write_bits_idx(MetadataArray_1_io_write_bits_idx),
    .io_write_bits_way_en(MetadataArray_1_io_write_bits_way_en),
    .io_write_bits_data_tag(MetadataArray_1_io_write_bits_data_tag),
    .io_write_bits_data_coh_state(MetadataArray_1_io_write_bits_data_coh_state),
    .io_resp_0_tag(MetadataArray_1_io_resp_0_tag),
    .io_resp_0_coh_state(MetadataArray_1_io_resp_0_coh_state)
  );
  AMOALU AMOALU_1 (
    .clk(AMOALU_1_clk),
    .reset(AMOALU_1_reset),
    .io_addr(AMOALU_1_io_addr),
    .io_cmd(AMOALU_1_io_cmd),
    .io_typ(AMOALU_1_io_typ),
    .io_lhs(AMOALU_1_io_lhs),
    .io_rhs(AMOALU_1_io_rhs),
    .io_out(AMOALU_1_io_out)
  );
  assign io_cpu_req_ready = GEN_13;
  assign io_cpu_s2_nack = GEN_115;
  assign io_cpu_resp_valid = GEN_111;
  assign io_cpu_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_cmd = s2_req_cmd;
  assign io_cpu_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_data = T_4493;
  assign io_cpu_resp_bits_replay = doUncachedResp;
  assign io_cpu_resp_bits_has_data = s2_read;
  assign io_cpu_resp_bits_data_word_bypass = T_4452;
  assign io_cpu_resp_bits_store_data = pstore1_data;
  assign io_cpu_replay_next = T_4419;
  assign io_cpu_xcpt_ma_ld = T_2884;
  assign io_cpu_xcpt_ma_st = T_2885;
  assign io_cpu_xcpt_pf_ld = T_2886;
  assign io_cpu_xcpt_pf_st = T_2887;
  assign io_cpu_ordered = T_4418;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_pum = tlb_io_ptw_req_bits_pum;
  assign io_ptw_req_bits_mxr = tlb_io_ptw_req_bits_mxr;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = T_3706;
  assign io_mem_acquire_bits_addr_block = GEN_63;
  assign io_mem_acquire_bits_client_xact_id = GEN_64;
  assign io_mem_acquire_bits_addr_beat = GEN_65;
  assign io_mem_acquire_bits_is_builtin_type = GEN_66;
  assign io_mem_acquire_bits_a_type = GEN_67;
  assign io_mem_acquire_bits_union = GEN_68;
  assign io_mem_acquire_bits_data = GEN_69;
  assign io_mem_probe_ready = T_3907;
  assign io_mem_release_valid = GEN_88;
  assign io_mem_release_bits_addr_beat = writebackCount;
  assign io_mem_release_bits_addr_block = probe_bits_addr_block;
  assign io_mem_release_bits_client_xact_id = GEN_101;
  assign io_mem_release_bits_voluntary = GEN_102;
  assign io_mem_release_bits_r_type = GEN_103;
  assign io_mem_release_bits_data = s2_data;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_finish_valid = fq_io_deq_valid;
  assign io_mem_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_3842;
  assign fq_io_enq_bits_manager_xact_id = T_3866_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_3866_manager_id;
  assign fq_io_deq_ready = io_mem_finish_ready;
  assign T_1924 = refillDone;
  assign T_1928 = T_1927[0];
  assign T_1929 = T_1927[2];
  assign T_1930 = T_1928 ^ T_1929;
  assign T_1931 = T_1927[3];
  assign T_1932 = T_1930 ^ T_1931;
  assign T_1933 = T_1927[5];
  assign T_1934 = T_1932 ^ T_1933;
  assign T_1935 = T_1927[15:1];
  assign T_1936 = {T_1934,T_1935};
  assign GEN_2 = T_1924 ? T_1936 : T_1927;
  assign metaReadArb_clk = clk;
  assign metaReadArb_reset = reset;
  assign metaReadArb_io_in_0_valid = flushing;
  assign metaReadArb_io_in_0_bits_idx = T_4517;
  assign metaReadArb_io_in_0_bits_way_en = 1'h1;
  assign metaReadArb_io_in_1_valid = T_3897;
  assign metaReadArb_io_in_1_bits_idx = io_mem_probe_bits_addr_block[5:0];
  assign metaReadArb_io_in_1_bits_way_en = 1'h1;
  assign metaReadArb_io_in_2_valid = io_cpu_req_valid;
  assign metaReadArb_io_in_2_bits_idx = T_2384;
  assign metaReadArb_io_in_2_bits_way_en = 1'h1;
  assign metaReadArb_io_out_ready = MetadataArray_1_io_read_ready;
  assign metaWriteArb_clk = clk;
  assign metaWriteArb_reset = reset;
  assign metaWriteArb_io_in_0_valid = T_3091;
  assign metaWriteArb_io_in_0_bits_idx = T_3092;
  assign metaWriteArb_io_in_0_bits_way_en = s2_victim_way[0];
  assign metaWriteArb_io_in_0_bits_data_tag = T_3160;
  assign metaWriteArb_io_in_0_bits_data_coh_state = T_3138_state;
  assign metaWriteArb_io_in_1_valid = refillDone;
  assign metaWriteArb_io_in_1_bits_idx = T_3092;
  assign metaWriteArb_io_in_1_bits_way_en = s2_victim_way[0];
  assign metaWriteArb_io_in_1_bits_data_tag = T_3160;
  assign metaWriteArb_io_in_1_bits_data_coh_state = T_3805_state;
  assign metaWriteArb_io_in_2_valid = T_4404;
  assign metaWriteArb_io_in_2_bits_idx = T_4408;
  assign metaWriteArb_io_in_2_bits_way_en = releaseWay[0];
  assign metaWriteArb_io_in_2_bits_data_tag = T_4412;
  assign metaWriteArb_io_in_2_bits_data_coh_state = newCoh_state;
  assign metaWriteArb_io_out_ready = MetadataArray_1_io_write_ready;
  assign data_clk = clk;
  assign data_reset = reset;
  assign data_io_req_valid = dataArb_io_out_valid;
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr;
  assign data_io_req_bits_write = dataArb_io_out_bits_write;
  assign data_io_req_bits_wdata = dataArb_io_out_bits_wdata;
  assign data_io_req_bits_wmask = dataArb_io_out_bits_wmask;
  assign data_io_req_bits_way_en = dataArb_io_out_bits_way_en;
  assign dataArb_clk = clk;
  assign dataArb_reset = reset;
  assign dataArb_io_in_0_valid = pstore_drain;
  assign dataArb_io_in_0_bits_addr = T_3031[11:0];
  assign dataArb_io_in_0_bits_write = 1'h1;
  assign dataArb_io_in_0_bits_wdata = T_3033;
  assign dataArb_io_in_0_bits_wmask = T_3077[7:0];
  assign dataArb_io_in_0_bits_way_en = T_3032;
  assign dataArb_io_in_1_valid = T_3753;
  assign dataArb_io_in_1_bits_addr = T_3764[11:0];
  assign dataArb_io_in_1_bits_write = 1'h1;
  assign dataArb_io_in_1_bits_wdata = io_mem_grant_bits_data;
  assign dataArb_io_in_1_bits_wmask = 8'hff;
  assign dataArb_io_in_1_bits_way_en = s2_victim_way[0];
  assign dataArb_io_in_2_valid = T_4395;
  assign dataArb_io_in_2_bits_addr = T_4399[11:0];
  assign dataArb_io_in_2_bits_write = 1'h0;
  assign dataArb_io_in_2_bits_wdata = GEN_14;
  assign dataArb_io_in_2_bits_wmask = GEN_31;
  assign dataArb_io_in_2_bits_way_en = 1'h1;
  assign dataArb_io_in_3_valid = T_2367;
  assign dataArb_io_in_3_bits_addr = io_cpu_req_bits_addr[11:0];
  assign dataArb_io_in_3_bits_write = 1'h0;
  assign dataArb_io_in_3_bits_wdata = GEN_32;
  assign dataArb_io_in_3_bits_wmask = GEN_77;
  assign dataArb_io_in_3_bits_way_en = 1'h1;
  assign dataArb_io_out_ready = 1'h1;
  assign T_2218 = io_cpu_req_ready & io_cpu_req_valid;
  assign T_2220 = io_mem_probe_ready & io_mem_probe_valid;
  assign GEN_3 = T_2220 ? io_mem_probe_bits_addr_block : probe_bits_addr_block;
  assign GEN_4 = T_2220 ? io_mem_probe_bits_p_type : probe_bits_p_type;
  assign s1_nack = GEN_109;
  assign T_2247 = io_cpu_s1_kill == 1'h0;
  assign T_2248 = s1_valid & T_2247;
  assign T_2249 = {io_cpu_xcpt_pf_ld,io_cpu_xcpt_pf_st};
  assign T_2250 = {io_cpu_xcpt_ma_ld,io_cpu_xcpt_ma_st};
  assign T_2251 = {T_2250,T_2249};
  assign T_2253 = T_2251 != 4'h0;
  assign T_2255 = T_2253 == 1'h0;
  assign s1_valid_masked = T_2248 & T_2255;
  assign T_2257 = s1_nack == 1'h0;
  assign s1_valid_not_nacked = s1_valid_masked & T_2257;
  assign T_2324 = io_cpu_req_bits_addr[39:12];
  assign T_2325 = io_cpu_req_bits_addr[5:0];
  assign T_2326 = {T_2324,metaReadArb_io_out_bits_idx};
  assign T_2327 = {T_2326,T_2325};
  assign GEN_5 = metaReadArb_io_out_valid ? T_2327 : s1_req_addr;
  assign GEN_6 = metaReadArb_io_out_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign GEN_7 = metaReadArb_io_out_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign GEN_8 = metaReadArb_io_out_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign GEN_9 = metaReadArb_io_out_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign GEN_10 = metaReadArb_io_out_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T_2328 = s1_req_cmd == 5'h0;
  assign T_2329 = s1_req_cmd == 5'h6;
  assign T_2330 = T_2328 | T_2329;
  assign T_2331 = s1_req_cmd == 5'h7;
  assign T_2332 = T_2330 | T_2331;
  assign T_2333 = s1_req_cmd[3];
  assign T_2334 = s1_req_cmd == 5'h4;
  assign T_2335 = T_2333 | T_2334;
  assign s1_read = T_2332 | T_2335;
  assign T_2336 = s1_req_cmd == 5'h1;
  assign T_2338 = T_2336 | T_2331;
  assign s1_write = T_2338 | T_2335;
  assign s1_readwrite = s1_read | s1_write;
  assign pstore1_valid = T_2979;
  assign T_2348 = release_state == 3'h2;
  assign T_2349 = release_state == 3'h3;
  assign inWriteback = T_2348 | T_2349;
  assign releaseWay = GEN_106;
  assign T_2351 = release_state == 3'h0;
  assign T_2353 = grant_wait == 1'h0;
  assign T_2354 = T_2351 & T_2353;
  assign T_2357 = T_2354 & T_2257;
  assign T_2358 = io_cpu_req_bits_cmd == 5'h0;
  assign T_2359 = io_cpu_req_bits_cmd == 5'h6;
  assign T_2360 = T_2358 | T_2359;
  assign T_2361 = io_cpu_req_bits_cmd == 5'h7;
  assign T_2362 = T_2360 | T_2361;
  assign T_2363 = io_cpu_req_bits_cmd[3];
  assign T_2364 = io_cpu_req_bits_cmd == 5'h4;
  assign T_2365 = T_2363 | T_2364;
  assign T_2366 = T_2362 | T_2365;
  assign T_2367 = io_cpu_req_valid & T_2366;
  assign T_2372 = dataArb_io_in_3_ready == 1'h0;
  assign T_2382 = T_2372 & T_2366;
  assign GEN_11 = T_2382 ? 1'h0 : T_2357;
  assign T_2384 = io_cpu_req_bits_addr[11:6];
  assign T_2388 = metaReadArb_io_in_2_ready == 1'h0;
  assign GEN_12 = T_2388 ? 1'h0 : GEN_11;
  assign tlb_clk = clk;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = T_2390;
  assign tlb_io_req_bits_vpn = T_2391;
  assign tlb_io_req_bits_passthrough = s1_req_phys;
  assign tlb_io_req_bits_instruction = 1'h0;
  assign tlb_io_req_bits_store = s1_write;
  assign tlb_io_ptw_req_ready = io_ptw_req_ready;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_hardware = io_ptw_resp_bits_pte_reserved_for_hardware;
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a;
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g;
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u;
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x;
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w;
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign tlb_io_ptw_ptbr_asid = io_ptw_ptbr_asid;
  assign tlb_io_ptw_ptbr_ppn = io_ptw_ptbr_ppn;
  assign tlb_io_ptw_invalidate = io_ptw_invalidate;
  assign tlb_io_ptw_status_debug = io_ptw_status_debug;
  assign tlb_io_ptw_status_prv = io_ptw_status_prv;
  assign tlb_io_ptw_status_sd = io_ptw_status_sd;
  assign tlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign tlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign tlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign tlb_io_ptw_status_vm = io_ptw_status_vm;
  assign tlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr;
  assign tlb_io_ptw_status_pum = io_ptw_status_pum;
  assign tlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign tlb_io_ptw_status_xs = io_ptw_status_xs;
  assign tlb_io_ptw_status_fs = io_ptw_status_fs;
  assign tlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign tlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign tlb_io_ptw_status_spp = io_ptw_status_spp;
  assign tlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign tlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign tlb_io_ptw_status_spie = io_ptw_status_spie;
  assign tlb_io_ptw_status_upie = io_ptw_status_upie;
  assign tlb_io_ptw_status_mie = io_ptw_status_mie;
  assign tlb_io_ptw_status_hie = io_ptw_status_hie;
  assign tlb_io_ptw_status_sie = io_ptw_status_sie;
  assign tlb_io_ptw_status_uie = io_ptw_status_uie;
  assign T_2390 = s1_valid_masked & s1_readwrite;
  assign T_2391 = s1_req_addr[39:12];
  assign T_2394 = tlb_io_req_ready == 1'h0;
  assign T_2396 = io_cpu_req_bits_phys == 1'h0;
  assign T_2397 = T_2394 & T_2396;
  assign GEN_13 = T_2397 ? 1'h0 : GEN_12;
  assign T_2399 = s1_valid & s1_readwrite;
  assign T_2400 = T_2399 & tlb_io_resp_miss;
  assign T_2402 = s1_req_addr[11:0];
  assign s1_paddr = {tlb_io_resp_ppn,T_2402};
  assign T_2403 = probe_bits_addr_block[25:6];
  assign T_2404 = s1_paddr[31:12];
  assign s1_tag = s1_probe ? T_2403 : T_2404;
  assign s1_victim_way = 1'h0;
  assign MetadataArray_1_clk = clk;
  assign MetadataArray_1_reset = reset;
  assign MetadataArray_1_io_read_valid = metaReadArb_io_out_valid;
  assign MetadataArray_1_io_read_bits_idx = metaReadArb_io_out_bits_idx;
  assign MetadataArray_1_io_read_bits_way_en = metaReadArb_io_out_bits_way_en;
  assign MetadataArray_1_io_write_valid = metaWriteArb_io_out_valid;
  assign MetadataArray_1_io_write_bits_idx = metaWriteArb_io_out_bits_idx;
  assign MetadataArray_1_io_write_bits_way_en = metaWriteArb_io_out_bits_way_en;
  assign MetadataArray_1_io_write_bits_data_tag = metaWriteArb_io_out_bits_data_tag;
  assign MetadataArray_1_io_write_bits_data_coh_state = metaWriteArb_io_out_bits_data_coh_state;
  assign T_2406 = MetadataArray_1_io_resp_0_coh_state != 2'h0;
  assign T_2407 = MetadataArray_1_io_resp_0_tag == s1_tag;
  assign s1_hit_way = T_2406 & T_2407;
  assign T_2431_state = 2'h0;
  assign T_2455 = T_2407 ? MetadataArray_1_io_resp_0_coh_state : 2'h0;
  assign s1_hit_state_state = T_2455;
  assign T_2587 = s1_probe | s2_probe;
  assign T_2588 = release_state != 3'h0;
  assign releaseInFlight = T_2587 | T_2588;
  assign s2_valid_masked = s2_valid & T_2591;
  assign T_2659 = s1_valid_not_nacked | s1_flush_valid;
  assign T_2661 = tlb_io_resp_cacheable == 1'h0;
  assign GEN_15 = T_2659 ? {{8'd0}, s1_paddr} : s2_req_addr;
  assign GEN_16 = T_2659 ? s1_req_tag : s2_req_tag;
  assign GEN_17 = T_2659 ? s1_req_cmd : s2_req_cmd;
  assign GEN_18 = T_2659 ? s1_req_typ : s2_req_typ;
  assign GEN_19 = T_2659 ? s1_req_phys : s2_req_phys;
  assign GEN_20 = T_2659 ? s1_req_data : s2_req_data;
  assign GEN_21 = T_2659 ? T_2661 : s2_uncached;
  assign T_2664 = s2_req_cmd == 5'h0;
  assign T_2665 = s2_req_cmd == 5'h6;
  assign T_2666 = T_2664 | T_2665;
  assign T_2667 = s2_req_cmd == 5'h7;
  assign T_2668 = T_2666 | T_2667;
  assign T_2669 = s2_req_cmd[3];
  assign T_2670 = s2_req_cmd == 5'h4;
  assign T_2671 = T_2669 | T_2670;
  assign s2_read = T_2668 | T_2671;
  assign T_2672 = s2_req_cmd == 5'h1;
  assign T_2674 = T_2672 | T_2667;
  assign s2_write = T_2674 | T_2671;
  assign s2_readwrite = s2_read | s2_write;
  assign T_2678 = s1_valid | inWriteback;
  assign GEN_22 = T_2678 ? data_io_resp_0 : s2_data;
  assign GEN_23 = s1_probe ? s1_hit_way : s2_probe_way;
  assign GEN_24 = s1_probe ? s1_hit_state_state : s2_probe_state_state;
  assign GEN_25 = s1_valid_not_nacked ? s1_hit_way : s2_hit_way;
  assign GEN_26 = s1_valid_not_nacked ? s1_hit_state_state : s2_hit_state_state;
  assign T_2728 = s2_req_cmd == 5'h3;
  assign T_2729 = s2_write | T_2728;
  assign T_2731 = T_2729 | T_2665;
  assign T_2732 = s2_hit_state_state == 2'h1;
  assign T_2733 = s2_hit_state_state == 2'h2;
  assign T_2734 = T_2732 | T_2733;
  assign s2_hit = T_2731 ? T_2734 : T_2734;
  assign T_2738 = s2_valid_masked & s2_readwrite;
  assign s2_valid_hit = T_2738 & s2_hit;
  assign T_2741 = s2_hit == 1'h0;
  assign T_2742 = T_2738 & T_2741;
  assign T_2743 = pstore1_valid | pstore2_valid;
  assign T_2745 = T_2743 == 1'h0;
  assign T_2746 = T_2742 & T_2745;
  assign T_2748 = release_ack_wait == 1'h0;
  assign s2_valid_miss = T_2746 & T_2748;
  assign T_2750 = s2_uncached == 1'h0;
  assign s2_valid_cached_miss = s2_valid_miss & T_2750;
  assign s2_victimize = s2_valid_cached_miss | s2_flush_valid;
  assign s2_valid_uncached = s2_valid_miss & s2_uncached;
  assign T_2751 = s2_hit_state_state != 2'h0;
  assign T_2753 = s2_flush_valid == 1'h0;
  assign T_2754 = T_2751 & T_2753;
  assign GEN_27 = T_2659 ? s1_victim_way : T_2756;
  assign T_2758 = 2'h1 << T_2756;
  assign s2_victim_way = T_2754 ? {{1'd0}, s2_hit_way} : T_2758;
  assign GEN_0_tag = GEN_28;
  assign GEN_0_coh_state = GEN_29;
  assign GEN_28 = MetadataArray_1_io_resp_0_tag;
  assign GEN_29 = MetadataArray_1_io_resp_0_coh_state;
  assign GEN_30 = T_2659 ? GEN_0_tag : s2_victim_tag;
  assign GEN_1_tag = GEN_28;
  assign GEN_1_coh_state = GEN_29;
  assign GEN_33 = T_2659 ? GEN_1_coh_state : T_2766_state;
  assign s2_victim_state_state = T_2754 ? s2_hit_state_state : T_2766_state;
  assign s2_victim_dirty = s2_victim_state_state == 2'h2;
  assign T_2816 = s2_write ? 2'h2 : s2_hit_state_state;
  assign s2_new_hit_state_state = T_2816;
  assign T_2860 = s2_hit_state_state == s2_new_hit_state_state;
  assign s2_update_meta = T_2860 == 1'h0;
  assign T_2863 = s2_valid_hit == 1'h0;
  assign T_2864 = s2_valid & T_2863;
  assign T_2865 = s2_valid_uncached & io_mem_acquire_ready;
  assign T_2867 = T_2865 == 1'h0;
  assign T_2868 = T_2864 & T_2867;
  assign T_2871 = T_2863 | s2_update_meta;
  assign T_2872 = s2_valid & T_2871;
  assign GEN_34 = T_2872 ? 1'h1 : T_2400;
  assign T_2875 = s1_req_typ[1:0];
  assign T_2877 = 4'h1 << T_2875;
  assign T_2879 = T_2877 - 4'h1;
  assign T_2880 = T_2879[3:0];
  assign T_2881 = T_2880[2:0];
  assign GEN_0 = {{37'd0}, T_2881};
  assign T_2882 = s1_req_addr & GEN_0;
  assign misaligned = T_2882 != 40'h0;
  assign T_2884 = s1_read & misaligned;
  assign T_2885 = s1_write & misaligned;
  assign T_2886 = s1_read & tlb_io_resp_xcpt_ld;
  assign T_2887 = s1_write & tlb_io_resp_xcpt_st;
  assign lrscValid = lrscCount > 5'h0;
  assign T_2895 = s2_req_addr[39:6];
  assign T_2896 = lrscAddr == T_2895;
  assign T_2897 = lrscValid & T_2896;
  assign T_2899 = T_2897 == 1'h0;
  assign s2_sc_fail = T_2667 & T_2899;
  assign T_2900 = s2_valid_hit & T_2665;
  assign GEN_35 = T_2900 ? 5'h1f : lrscCount;
  assign GEN_36 = T_2900 ? T_2895 : lrscAddr;
  assign T_2904 = lrscCount - 5'h1;
  assign T_2905 = T_2904[4:0];
  assign GEN_37 = lrscValid ? T_2905 : GEN_35;
  assign T_2906 = s2_valid_hit & T_2667;
  assign T_2907 = T_2906 | io_cpu_invalidate_lr;
  assign GEN_38 = T_2907 ? 5'h0 : GEN_37;
  assign T_2909 = s1_valid_not_nacked & s1_write;
  assign GEN_39 = T_2909 ? s1_req_cmd : pstore1_cmd;
  assign GEN_40 = T_2909 ? s1_req_typ : pstore1_typ;
  assign GEN_41 = T_2909 ? s1_paddr : pstore1_addr;
  assign GEN_42 = T_2909 ? io_cpu_s1_data : pstore1_data;
  assign GEN_43 = T_2909 ? s1_hit_way : pstore1_way;
  assign T_2914 = pstore1_typ[1:0];
  assign T_2916 = T_2914 == 2'h0;
  assign T_2917 = pstore1_data[7:0];
  assign T_2918 = {T_2917,T_2917};
  assign T_2919 = {T_2918,T_2918};
  assign T_2920 = {T_2919,T_2919};
  assign T_2922 = T_2914 == 2'h1;
  assign T_2923 = pstore1_data[15:0];
  assign T_2924 = {T_2923,T_2923};
  assign T_2925 = {T_2924,T_2924};
  assign T_2927 = T_2914 == 2'h2;
  assign T_2928 = pstore1_data[31:0];
  assign T_2929 = {T_2928,T_2928};
  assign T_2930 = T_2927 ? T_2929 : pstore1_data;
  assign T_2931 = T_2922 ? T_2925 : T_2930;
  assign T_2932 = T_2916 ? T_2920 : T_2931;
  assign pstore1_storegen_data = AMOALU_1_io_out;
  assign T_2934 = pstore1_cmd == 5'h0;
  assign T_2935 = pstore1_cmd == 5'h6;
  assign T_2936 = T_2934 | T_2935;
  assign T_2937 = pstore1_cmd == 5'h7;
  assign T_2938 = T_2936 | T_2937;
  assign T_2939 = pstore1_cmd[3];
  assign T_2940 = pstore1_cmd == 5'h4;
  assign T_2941 = T_2939 | T_2940;
  assign T_2942 = T_2938 | T_2941;
  assign T_2943 = pstore1_valid & pstore2_valid;
  assign T_2944 = s1_valid & s1_write;
  assign T_2945 = T_2944 | T_2942;
  assign pstore_drain_structural = T_2943 & T_2945;
  assign pstore_drain_opportunistic = T_2367 == 1'h0;
  assign pstore_drain_on_miss = releaseInFlight | io_cpu_s2_nack;
  assign T_2960 = T_2942 == 1'h0;
  assign T_2961 = pstore1_valid & T_2960;
  assign T_2962 = T_2961 | pstore2_valid;
  assign T_2963 = pstore_drain_opportunistic | pstore_drain_on_miss;
  assign T_2964 = T_2962 & T_2963;
  assign pstore_drain = pstore_drain_structural | T_2964;
  assign T_2965 = s2_valid_hit & s2_write;
  assign T_2967 = s2_sc_fail == 1'h0;
  assign T_2968 = T_2965 & T_2967;
  assign T_2972 = T_2968 == 1'h0;
  assign T_2974 = T_2970 == 1'h0;
  assign T_2975 = T_2972 | T_2974;
  assign T_2976 = T_2975 | reset;
  assign T_2978 = T_2976 == 1'h0;
  assign T_2979 = T_2968 | T_2970;
  assign T_2980 = T_2979 & pstore2_valid;
  assign T_2982 = pstore_drain == 1'h0;
  assign T_2983 = T_2980 & T_2982;
  assign T_2985 = pstore2_valid == pstore_drain;
  assign advance_pstore1 = pstore1_valid & T_2985;
  assign T_2988 = pstore2_valid & T_2982;
  assign T_2989 = T_2988 | advance_pstore1;
  assign GEN_44 = advance_pstore1 ? pstore1_addr : pstore2_addr;
  assign GEN_45 = advance_pstore1 ? pstore1_way : pstore2_way;
  assign GEN_46 = advance_pstore1 ? pstore1_storegen_data : pstore2_storegen_data;
  assign T_2991 = pstore1_addr[0];
  assign T_2995 = T_2914 >= 2'h1;
  assign T_2999 = T_2991 | T_2995;
  assign T_3002 = T_2991 ? 1'h0 : 1'h1;
  assign T_3003 = {T_2999,T_3002};
  assign T_3004 = pstore1_addr[1];
  assign T_3006 = T_3004 ? T_3003 : 2'h0;
  assign T_3008 = T_2914 >= 2'h2;
  assign T_3011 = T_3008 ? 2'h3 : 2'h0;
  assign T_3012 = T_3006 | T_3011;
  assign T_3015 = T_3004 ? 2'h0 : T_3003;
  assign T_3016 = {T_3012,T_3015};
  assign T_3017 = pstore1_addr[2];
  assign T_3019 = T_3017 ? T_3016 : 4'h0;
  assign T_3021 = T_2914 >= 2'h3;
  assign T_3024 = T_3021 ? 4'hf : 4'h0;
  assign T_3025 = T_3019 | T_3024;
  assign T_3028 = T_3017 ? 4'h0 : T_3016;
  assign T_3029 = {T_3025,T_3028};
  assign GEN_47 = advance_pstore1 ? T_3029 : pstore2_storegen_mask;
  assign T_3031 = pstore2_valid ? pstore2_addr : pstore1_addr;
  assign T_3032 = pstore2_valid ? pstore2_way : pstore1_way;
  assign T_3033 = pstore2_valid ? pstore2_storegen_data : pstore1_storegen_data;
  assign T_3076 = pstore2_valid ? pstore2_storegen_mask : T_3029;
  assign GEN_1 = {{15'd0}, T_3076};
  assign T_3077 = GEN_1 << 4'h0;
  assign s1_idx = s1_req_addr[11:3];
  assign T_3078 = pstore1_addr[11:3];
  assign T_3079 = T_3078 == s1_idx;
  assign T_3080 = pstore1_valid & T_3079;
  assign T_3081 = pstore2_addr[11:3];
  assign T_3082 = T_3081 == s1_idx;
  assign T_3083 = pstore2_valid & T_3082;
  assign T_3084 = T_3080 | T_3083;
  assign s1_raw_hazard = s1_read & T_3084;
  assign T_3085 = s1_valid & s1_raw_hazard;
  assign GEN_48 = T_3085 ? 1'h1 : GEN_34;
  assign T_3087 = s2_valid_hit & s2_update_meta;
  assign T_3089 = s2_victim_dirty == 1'h0;
  assign T_3090 = s2_victimize & T_3089;
  assign T_3091 = T_3087 | T_3090;
  assign T_3092 = s2_req_addr[11:6];
  assign T_3116_state = 2'h0;
  assign T_3138_state = s2_valid_hit ? s2_new_hit_state_state : T_3116_state;
  assign T_3160 = s2_req_addr[31:12];
  assign T_3162 = s2_req_addr[31:6];
  assign T_3177 = {s2_req_cmd,1'h1};
  assign cachedGetMessage_addr_block = T_3162;
  assign cachedGetMessage_client_xact_id = 1'h0;
  assign cachedGetMessage_addr_beat = 3'h0;
  assign cachedGetMessage_is_builtin_type = 1'h0;
  assign cachedGetMessage_a_type = {{2'd0}, T_2731};
  assign cachedGetMessage_union = {{5'd0}, T_3177};
  assign cachedGetMessage_data = 64'h0;
  assign T_3237 = s2_req_addr[5:3];
  assign T_3238 = s2_req_addr[2:0];
  assign T_3269 = s2_req_typ[1:0];
  assign T_3279 = {T_3238,T_3269};
  assign T_3280 = {T_3279,6'h0};
  assign uncachedGetMessage_addr_block = T_3162;
  assign uncachedGetMessage_client_xact_id = 1'h0;
  assign uncachedGetMessage_addr_beat = T_3237;
  assign uncachedGetMessage_is_builtin_type = 1'h1;
  assign uncachedGetMessage_a_type = 3'h0;
  assign uncachedGetMessage_union = T_3280;
  assign uncachedGetMessage_data = 64'h0;
  assign GEN_125 = {{15'd0}, T_3029};
  assign T_3427 = GEN_125 << 4'h0;
  assign T_3465 = T_3427[7:0];
  assign T_3475 = {T_3465,1'h0};
  assign T_3495 = {{2'd0}, T_3475};
  assign uncachedPutMessage_addr_block = T_3162;
  assign uncachedPutMessage_client_xact_id = 1'h0;
  assign uncachedPutMessage_addr_beat = T_3237;
  assign uncachedPutMessage_is_builtin_type = 1'h1;
  assign uncachedPutMessage_a_type = 3'h2;
  assign uncachedPutMessage_union = T_3495;
  assign uncachedPutMessage_data = T_2932;
  assign T_3617 = {T_3279,T_3177};
  assign uncachedPutAtomicMessage_addr_block = T_3162;
  assign uncachedPutAtomicMessage_client_xact_id = 1'h0;
  assign uncachedPutAtomicMessage_addr_beat = T_3237;
  assign uncachedPutAtomicMessage_is_builtin_type = 1'h1;
  assign uncachedPutAtomicMessage_a_type = 3'h4;
  assign uncachedPutAtomicMessage_union = T_3617;
  assign uncachedPutAtomicMessage_data = T_2932;
  assign T_3704 = s2_valid_cached_miss & T_3089;
  assign T_3705 = T_3704 | s2_valid_uncached;
  assign T_3706 = T_3705 & fq_io_enq_ready;
  assign T_3708 = s2_valid_masked == 1'h0;
  assign T_3711 = T_2751 == 1'h0;
  assign T_3712 = T_3708 | T_3711;
  assign T_3713 = T_3712 | reset;
  assign T_3715 = T_3713 == 1'h0;
  assign GEN_49 = T_2942 ? uncachedPutAtomicMessage_addr_block : uncachedPutMessage_addr_block;
  assign GEN_50 = T_2942 ? uncachedPutAtomicMessage_client_xact_id : uncachedPutMessage_client_xact_id;
  assign GEN_51 = T_2942 ? uncachedPutAtomicMessage_addr_beat : uncachedPutMessage_addr_beat;
  assign GEN_52 = T_2942 ? uncachedPutAtomicMessage_is_builtin_type : uncachedPutMessage_is_builtin_type;
  assign GEN_53 = T_2942 ? uncachedPutAtomicMessage_a_type : uncachedPutMessage_a_type;
  assign GEN_54 = T_2942 ? uncachedPutAtomicMessage_union : uncachedPutMessage_union;
  assign GEN_55 = T_2942 ? uncachedPutAtomicMessage_data : uncachedPutMessage_data;
  assign GEN_56 = s2_write ? GEN_49 : uncachedGetMessage_addr_block;
  assign GEN_57 = s2_write ? GEN_50 : uncachedGetMessage_client_xact_id;
  assign GEN_58 = s2_write ? GEN_51 : uncachedGetMessage_addr_beat;
  assign GEN_59 = s2_write ? GEN_52 : uncachedGetMessage_is_builtin_type;
  assign GEN_60 = s2_write ? GEN_53 : uncachedGetMessage_a_type;
  assign GEN_61 = s2_write ? GEN_54 : uncachedGetMessage_union;
  assign GEN_62 = s2_write ? GEN_55 : uncachedGetMessage_data;
  assign GEN_63 = s2_uncached ? GEN_56 : cachedGetMessage_addr_block;
  assign GEN_64 = s2_uncached ? GEN_57 : cachedGetMessage_client_xact_id;
  assign GEN_65 = s2_uncached ? GEN_58 : cachedGetMessage_addr_beat;
  assign GEN_66 = s2_uncached ? GEN_59 : cachedGetMessage_is_builtin_type;
  assign GEN_67 = s2_uncached ? GEN_60 : cachedGetMessage_a_type;
  assign GEN_68 = s2_uncached ? GEN_61 : cachedGetMessage_union;
  assign GEN_69 = s2_uncached ? GEN_62 : cachedGetMessage_data;
  assign T_3716 = io_mem_acquire_ready & io_mem_acquire_valid;
  assign GEN_70 = T_3716 ? 1'h1 : grant_wait;
  assign T_3725_0 = 3'h5;
  assign GEN_126 = {{1'd0}, T_3725_0};
  assign T_3727 = io_mem_grant_bits_g_type == GEN_126;
  assign T_3728 = io_mem_grant_bits_g_type == 4'h0;
  assign T_3729 = io_mem_grant_bits_is_builtin_type ? T_3727 : T_3728;
  assign grantIsVoluntary = io_mem_grant_bits_is_builtin_type & T_3728;
  assign T_3733 = T_3729 == 1'h0;
  assign T_3735 = grantIsVoluntary == 1'h0;
  assign grantIsUncached = T_3733 & T_3735;
  assign T_3736 = grantIsVoluntary & release_ack_wait;
  assign T_3737 = grant_wait | T_3736;
  assign T_3738 = T_3737 | reset;
  assign T_3740 = T_3738 == 1'h0;
  assign GEN_71 = grantIsUncached ? io_mem_grant_bits_data : GEN_22;
  assign GEN_72 = grantIsVoluntary ? 1'h0 : release_ack_wait;
  assign GEN_73 = io_mem_grant_valid ? GEN_71 : GEN_22;
  assign GEN_74 = io_mem_grant_valid ? GEN_72 : release_ack_wait;
  assign T_3742 = io_mem_grant_ready & io_mem_grant_valid;
  assign T_3743 = T_3742 & T_3729;
  assign T_3746 = refillCount == 3'h7;
  assign T_3748 = refillCount + 3'h1;
  assign T_3749 = T_3748[2:0];
  assign GEN_75 = T_3743 ? T_3749 : refillCount;
  assign refillDone = T_3743 & T_3746;
  assign grantDone = refillDone | grantIsUncached;
  assign T_3751 = T_3742 & grantDone;
  assign GEN_76 = T_3751 ? 1'h0 : GEN_70;
  assign T_3753 = T_3729 & io_mem_grant_valid;
  assign T_3756 = dataArb_io_in_1_valid == 1'h0;
  assign T_3757 = dataArb_io_in_1_ready | T_3756;
  assign T_3758 = T_3757 | reset;
  assign T_3760 = T_3758 == 1'h0;
  assign T_3763 = {T_3162,io_mem_grant_bits_addr_beat};
  assign GEN_127 = {{3'd0}, T_3763};
  assign T_3764 = GEN_127 << 3;
  assign T_3768 = metaWriteArb_io_in_1_valid == 1'h0;
  assign T_3769 = T_3768 | metaWriteArb_io_in_1_ready;
  assign T_3770 = T_3769 | reset;
  assign T_3772 = T_3770 == 1'h0;
  assign T_3781 = s2_write ? 2'h2 : 2'h1;
  assign T_3782 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T_3781;
  assign T_3805_state = T_3782;
  assign T_3838 = T_3742 & T_3735;
  assign T_3841 = T_3733 | refillDone;
  assign T_3842 = T_3838 & T_3841;
  assign T_3866_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign T_3866_manager_id = io_mem_grant_bits_manager_id;
  assign T_3889 = fq_io_enq_ready | reset;
  assign T_3891 = T_3889 == 1'h0;
  assign T_3893 = releaseInFlight | lrscValid;
  assign block_probe = T_3893 | T_2900;
  assign T_3896 = block_probe == 1'h0;
  assign T_3897 = io_mem_probe_valid & T_3896;
  assign T_3900 = metaReadArb_io_in_1_ready & T_3896;
  assign T_3902 = s1_valid == 1'h0;
  assign T_3903 = T_3900 & T_3902;
  assign T_3905 = s2_valid == 1'h0;
  assign T_3906 = T_3905 | s2_valid_hit;
  assign T_3907 = T_3903 & T_3906;
  assign T_3910 = io_mem_release_ready & io_mem_release_valid;
  assign T_3911 = T_3910 & inWriteback;
  assign T_3914 = writebackCount == 3'h7;
  assign T_3916 = writebackCount + 3'h1;
  assign T_3917 = T_3916[2:0];
  assign GEN_78 = T_3911 ? T_3917 : writebackCount;
  assign writebackDone = T_3911 & T_3914;
  assign T_3920 = inWriteback == 1'h0;
  assign T_3921 = T_3910 & T_3920;
  assign releaseDone = writebackDone | T_3921;
  assign T_3923 = io_mem_release_ready == 1'h0;
  assign releaseRejected = io_mem_release_valid & T_3923;
  assign T_3924 = dataArb_io_in_2_ready & dataArb_io_in_2_valid;
  assign T_3926 = releaseRejected == 1'h0;
  assign T_3927 = s1_release_data_valid & T_3926;
  assign T_3929 = {1'h0,writebackCount};
  assign T_3932 = {1'h0,s2_release_data_valid};
  assign GEN_128 = {{1'd0}, s1_release_data_valid};
  assign T_3933 = GEN_128 + T_3932;
  assign T_3934 = T_3933[1:0];
  assign T_3935 = releaseRejected ? 2'h0 : T_3934;
  assign GEN_129 = {{2'd0}, T_3935};
  assign T_3936 = T_3929 + GEN_129;
  assign releaseDataBeat = T_3936[3:0];
  assign T_3960_state = 2'h0;
  assign T_3985 = T_3960_state == 2'h2;
  assign T_3986 = T_3985 ? 3'h0 : 3'h3;
  assign T_4015 = 2'h2 == probe_bits_p_type;
  assign T_4016 = T_4015 ? T_3986 : 3'h3;
  assign T_4017 = 2'h1 == probe_bits_p_type;
  assign T_4018 = T_4017 ? T_3986 : T_4016;
  assign T_4019 = 2'h0 == probe_bits_p_type;
  assign T_4020 = T_4019 ? T_3986 : T_4018;
  assign T_4049_addr_beat = 3'h0;
  assign T_4049_addr_block = probe_bits_addr_block;
  assign T_4049_client_xact_id = 1'h0;
  assign T_4049_voluntary = 1'h0;
  assign T_4049_r_type = T_4020;
  assign T_4049_data = 64'h0;
  assign T_4082 = s2_victim_dirty ? 3'h0 : 3'h3;
  assign voluntaryReleaseMessage_addr_beat = 3'h0;
  assign voluntaryReleaseMessage_addr_block = 26'h0;
  assign voluntaryReleaseMessage_client_xact_id = 1'h0;
  assign voluntaryReleaseMessage_voluntary = 1'h1;
  assign voluntaryReleaseMessage_r_type = T_4082;
  assign voluntaryReleaseMessage_data = 64'h0;
  assign voluntaryNewCoh_state = 2'h0;
  assign T_4196 = s2_probe_state_state == 2'h2;
  assign T_4197 = T_4196 ? 3'h0 : 3'h3;
  assign T_4227 = T_4015 ? T_4197 : 3'h3;
  assign T_4229 = T_4017 ? T_4197 : T_4227;
  assign T_4231 = T_4019 ? T_4197 : T_4229;
  assign probeResponseMessage_addr_beat = 3'h0;
  assign probeResponseMessage_addr_block = probe_bits_addr_block;
  assign probeResponseMessage_client_xact_id = 1'h0;
  assign probeResponseMessage_voluntary = 1'h0;
  assign probeResponseMessage_r_type = T_4231;
  assign probeResponseMessage_data = 64'h0;
  assign T_4287 = T_4015 ? 2'h0 : s2_probe_state_state;
  assign T_4289 = T_4017 ? 2'h0 : T_4287;
  assign T_4291 = T_4019 ? 2'h0 : T_4289;
  assign probeNewCoh_state = T_4291;
  assign newCoh_state = GEN_105;
  assign T_4356 = s2_victimize & s2_victim_dirty;
  assign T_4358 = s2_valid & T_2751;
  assign T_4360 = T_4358 == 1'h0;
  assign T_4361 = T_4360 | reset;
  assign T_4363 = T_4361 == 1'h0;
  assign T_4365 = {s2_victim_tag,T_3092};
  assign GEN_79 = T_4356 ? 3'h2 : release_state;
  assign GEN_80 = T_4356 ? T_4365 : GEN_3;
  assign GEN_81 = T_4196 ? 3'h3 : GEN_79;
  assign T_4367 = s2_probe_state_state != 2'h0;
  assign T_4369 = T_4196 == 1'h0;
  assign T_4370 = T_4369 & T_4367;
  assign GEN_82 = T_4370 ? 3'h4 : GEN_81;
  assign T_4374 = T_4367 == 1'h0;
  assign T_4375 = T_4369 & T_4374;
  assign GEN_83 = T_4375 ? 1'h1 : s2_release_data_valid;
  assign GEN_84 = T_4375 ? 3'h5 : GEN_82;
  assign GEN_85 = s2_probe ? GEN_84 : GEN_79;
  assign GEN_86 = s2_probe ? GEN_83 : s2_release_data_valid;
  assign GEN_87 = releaseDone ? 3'h0 : GEN_85;
  assign T_4377 = release_state == 3'h5;
  assign T_4378 = release_state == 3'h4;
  assign T_4379 = T_4377 | T_4378;
  assign GEN_88 = T_4379 ? 1'h1 : GEN_86;
  assign T_4383 = T_4378 | T_2349;
  assign GEN_89 = releaseDone ? 3'h7 : GEN_87;
  assign GEN_92 = T_4383 ? probeResponseMessage_client_xact_id : T_4049_client_xact_id;
  assign GEN_93 = T_4383 ? probeResponseMessage_voluntary : T_4049_voluntary;
  assign GEN_94 = T_4383 ? probeResponseMessage_r_type : T_4049_r_type;
  assign GEN_96 = T_4383 ? GEN_89 : GEN_87;
  assign T_4385 = release_state == 3'h6;
  assign T_4386 = T_2348 | T_4385;
  assign GEN_97 = releaseDone ? 3'h6 : GEN_96;
  assign GEN_98 = releaseDone ? 1'h1 : GEN_74;
  assign GEN_101 = T_4386 ? voluntaryReleaseMessage_client_xact_id : GEN_92;
  assign GEN_102 = T_4386 ? voluntaryReleaseMessage_voluntary : GEN_93;
  assign GEN_103 = T_4386 ? voluntaryReleaseMessage_r_type : GEN_94;
  assign GEN_105 = T_4386 ? voluntaryNewCoh_state : probeNewCoh_state;
  assign GEN_106 = T_4386 ? s2_victim_way : {{1'd0}, s2_probe_way};
  assign GEN_107 = T_4386 ? GEN_97 : GEN_96;
  assign GEN_108 = T_4386 ? GEN_98 : GEN_74;
  assign T_4390 = T_3910 == 1'h0;
  assign T_4391 = s2_probe & T_4390;
  assign GEN_109 = T_4391 ? 1'h1 : GEN_48;
  assign T_4394 = releaseDataBeat < 4'h8;
  assign T_4395 = inWriteback & T_4394;
  assign T_4397 = releaseDataBeat[2:0];
  assign T_4398 = {io_mem_release_bits_addr_block,T_4397};
  assign GEN_130 = {{3'd0}, T_4398};
  assign T_4399 = GEN_130 << 3;
  assign T_4403 = release_state == 3'h7;
  assign T_4404 = T_4385 | T_4403;
  assign T_4406 = {io_mem_release_bits_addr_block,io_mem_release_bits_addr_beat};
  assign T_4407 = {T_4406,3'h0};
  assign T_4408 = T_4407[11:6];
  assign T_4412 = T_4407[31:12];
  assign T_4413 = metaWriteArb_io_in_2_ready & metaWriteArb_io_in_2_valid;
  assign GEN_110 = T_4413 ? 3'h0 : GEN_107;
  assign T_4415 = s1_valid | s2_valid;
  assign T_4416 = T_4415 | grant_wait;
  assign T_4418 = T_4416 == 1'h0;
  assign T_4419 = io_mem_grant_valid & grantIsUncached;
  assign T_4422 = T_2863 | reset;
  assign T_4424 = T_4422 == 1'h0;
  assign GEN_111 = doUncachedResp ? 1'h1 : s2_valid_hit;
  assign s2_data_word = s2_data >> 7'h0;
  assign T_4429 = s2_req_typ[2];
  assign T_4431 = T_4429 == 1'h0;
  assign T_4433 = s2_req_addr[2];
  assign T_4434 = s2_data_word[63:32];
  assign T_4435 = s2_data_word[31:0];
  assign T_4436 = T_4433 ? T_4434 : T_4435;
  assign T_4442 = T_3269 == 2'h2;
  assign T_4444 = T_4436[31];
  assign T_4445 = T_4431 & T_4444;
  assign T_4449 = T_4445 ? 32'hffffffff : 32'h0;
  assign T_4451 = T_4442 ? T_4449 : T_4434;
  assign T_4452 = {T_4451,T_4436};
  assign T_4453 = s2_req_addr[1];
  assign T_4454 = T_4452[31:16];
  assign T_4455 = T_4452[15:0];
  assign T_4456 = T_4453 ? T_4454 : T_4455;
  assign T_4462 = T_3269 == 2'h1;
  assign T_4464 = T_4456[15];
  assign T_4465 = T_4431 & T_4464;
  assign T_4469 = T_4465 ? 48'hffffffffffff : 48'h0;
  assign T_4470 = T_4452[63:16];
  assign T_4471 = T_4462 ? T_4469 : T_4470;
  assign T_4472 = {T_4471,T_4456};
  assign T_4473 = s2_req_addr[0];
  assign T_4474 = T_4472[15:8];
  assign T_4475 = T_4472[7:0];
  assign T_4476 = T_4473 ? T_4474 : T_4475;
  assign T_4480 = T_2667 ? 8'h0 : T_4476;
  assign T_4482 = T_3269 == 2'h0;
  assign T_4483 = T_4482 | T_2667;
  assign T_4484 = T_4480[7];
  assign T_4485 = T_4431 & T_4484;
  assign T_4489 = T_4485 ? 56'hffffffffffffff : 56'h0;
  assign T_4490 = T_4472[63:8];
  assign T_4491 = T_4483 ? T_4489 : T_4490;
  assign T_4492 = {T_4491,T_4480};
  assign GEN_131 = {{63'd0}, s2_sc_fail};
  assign T_4493 = T_4492 | GEN_131;
  assign AMOALU_1_clk = clk;
  assign AMOALU_1_reset = reset;
  assign AMOALU_1_io_addr = pstore1_addr[2:0];
  assign AMOALU_1_io_cmd = pstore1_cmd;
  assign AMOALU_1_io_typ = pstore1_typ[1:0];
  assign AMOALU_1_io_lhs = s2_data_word;
  assign AMOALU_1_io_rhs = pstore1_data;
  assign T_4521 = T_3716 & T_2750;
  assign GEN_113 = T_4521 ? 1'h0 : flushed;
  assign T_4523 = s2_req_cmd == 5'h5;
  assign T_4524 = s2_valid_masked & T_4523;
  assign T_4526 = flushed == 1'h0;
  assign GEN_114 = T_4526 ? T_2748 : flushing;
  assign GEN_115 = T_4524 ? T_4526 : T_2868;
  assign GEN_116 = T_4524 ? GEN_114 : flushing;
  assign T_4531 = metaReadArb_io_in_0_ready & metaReadArb_io_in_0_valid;
  assign T_4533 = s1_flush_valid == 1'h0;
  assign T_4534 = T_4531 & T_4533;
  assign T_4537 = T_4534 & T_2753;
  assign T_4539 = T_4537 & T_2351;
  assign T_4542 = T_4539 & T_2748;
  assign T_4547 = T_4517 == 6'h3f;
  assign T_4549 = T_4517 + 6'h1;
  assign T_4550 = T_4549[5:0];
  assign GEN_117 = T_4547 ? 1'h1 : GEN_113;
  assign GEN_118 = s2_flush_valid ? T_4550 : T_4517;
  assign GEN_119 = s2_flush_valid ? GEN_117 : GEN_113;
  assign T_4553 = flushed & T_2351;
  assign T_4556 = T_4553 & T_2748;
  assign GEN_120 = T_4556 ? 1'h0 : GEN_116;
  assign GEN_122 = flushing ? GEN_118 : T_4517;
  assign GEN_123 = flushing ? GEN_119 : GEN_113;
  assign GEN_124 = flushing ? GEN_120 : GEN_116;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_14 = GEN_179[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_180[7:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_32 = GEN_181[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_77 = GEN_182[7:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {1{$random}};
  T_1927 = GEN_90[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {1{$random}};
  s1_valid = GEN_91[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_95 = {1{$random}};
  s1_probe = GEN_95[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_99 = {1{$random}};
  probe_bits_addr_block = GEN_99[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {1{$random}};
  probe_bits_p_type = GEN_100[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_104 = {2{$random}};
  s1_req_addr = GEN_104[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {1{$random}};
  s1_req_tag = GEN_112[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_121 = {1{$random}};
  s1_req_cmd = GEN_121[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_132 = {1{$random}};
  s1_req_typ = GEN_132[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_133 = {1{$random}};
  s1_req_phys = GEN_133[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_134 = {2{$random}};
  s1_req_data = GEN_134[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_135 = {1{$random}};
  s1_flush_valid = GEN_135[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_136 = {1{$random}};
  grant_wait = GEN_136[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_137 = {1{$random}};
  release_ack_wait = GEN_137[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_138 = {1{$random}};
  release_state = GEN_138[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_139 = {1{$random}};
  pstore2_valid = GEN_139[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_140 = {1{$random}};
  s2_valid = GEN_140[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_141 = {1{$random}};
  s2_probe = GEN_141[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_142 = {1{$random}};
  T_2591 = GEN_142[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_143 = {2{$random}};
  s2_req_addr = GEN_143[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_144 = {1{$random}};
  s2_req_tag = GEN_144[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_145 = {1{$random}};
  s2_req_cmd = GEN_145[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_146 = {1{$random}};
  s2_req_typ = GEN_146[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_147 = {1{$random}};
  s2_req_phys = GEN_147[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_148 = {2{$random}};
  s2_req_data = GEN_148[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_149 = {1{$random}};
  s2_uncached = GEN_149[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_150 = {1{$random}};
  s2_flush_valid = GEN_150[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_151 = {2{$random}};
  s2_data = GEN_151[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_152 = {1{$random}};
  s2_probe_way = GEN_152[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_153 = {1{$random}};
  s2_probe_state_state = GEN_153[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_154 = {1{$random}};
  s2_hit_way = GEN_154[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_155 = {1{$random}};
  s2_hit_state_state = GEN_155[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_156 = {1{$random}};
  T_2756 = GEN_156[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_157 = {1{$random}};
  s2_victim_tag = GEN_157[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_158 = {1{$random}};
  T_2766_state = GEN_158[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_159 = {1{$random}};
  lrscCount = GEN_159[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_160 = {2{$random}};
  lrscAddr = GEN_160[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_161 = {1{$random}};
  pstore1_cmd = GEN_161[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_162 = {1{$random}};
  pstore1_typ = GEN_162[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_163 = {1{$random}};
  pstore1_addr = GEN_163[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_164 = {2{$random}};
  pstore1_data = GEN_164[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_165 = {1{$random}};
  pstore1_way = GEN_165[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_166 = {1{$random}};
  T_2970 = GEN_166[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_167 = {1{$random}};
  pstore2_addr = GEN_167[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_168 = {1{$random}};
  pstore2_way = GEN_168[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_169 = {2{$random}};
  pstore2_storegen_data = GEN_169[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_170 = {1{$random}};
  pstore2_storegen_mask = GEN_170[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_171 = {1{$random}};
  refillCount = GEN_171[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_172 = {1{$random}};
  writebackCount = GEN_172[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_173 = {1{$random}};
  s1_release_data_valid = GEN_173[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_174 = {1{$random}};
  s2_release_data_valid = GEN_174[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_175 = {1{$random}};
  doUncachedResp = GEN_175[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_176 = {1{$random}};
  flushed = GEN_176[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_177 = {1{$random}};
  flushing = GEN_177[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_178 = {1{$random}};
  T_4517 = GEN_178[5:0];
  `endif
  GEN_179 = {2{$random}};
  GEN_180 = {1{$random}};
  GEN_181 = {2{$random}};
  GEN_182 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1927 <= 16'h1;
    end else begin
      if(T_1924) begin
        T_1927 <= T_1936;
      end
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_2218;
    end
    if(reset) begin
      s1_probe <= 1'h0;
    end else begin
      s1_probe <= T_2220;
    end
    if(1'h0) begin
    end else begin
      if(T_4356) begin
        probe_bits_addr_block <= T_4365;
      end else begin
        if(T_2220) begin
          probe_bits_addr_block <= io_mem_probe_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2220) begin
        probe_bits_p_type <= io_mem_probe_bits_p_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_addr <= T_2327;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_tag <= io_cpu_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_cmd <= io_cpu_req_bits_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_typ <= io_cpu_req_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_phys <= io_cpu_req_bits_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_data <= io_cpu_req_bits_data;
      end
    end
    if(1'h0) begin
    end else begin
      s1_flush_valid <= T_4542;
    end
    if(reset) begin
      grant_wait <= 1'h0;
    end else begin
      if(T_3751) begin
        grant_wait <= 1'h0;
      end else begin
        if(T_3716) begin
          grant_wait <= 1'h1;
        end
      end
    end
    if(reset) begin
      release_ack_wait <= 1'h0;
    end else begin
      if(T_4386) begin
        if(releaseDone) begin
          release_ack_wait <= 1'h1;
        end else begin
          if(io_mem_grant_valid) begin
            if(grantIsVoluntary) begin
              release_ack_wait <= 1'h0;
            end
          end
        end
      end else begin
        if(io_mem_grant_valid) begin
          if(grantIsVoluntary) begin
            release_ack_wait <= 1'h0;
          end
        end
      end
    end
    if(reset) begin
      release_state <= 3'h0;
    end else begin
      if(T_4413) begin
        release_state <= 3'h0;
      end else begin
        if(T_4386) begin
          if(releaseDone) begin
            release_state <= 3'h6;
          end else begin
            if(T_4383) begin
              if(releaseDone) begin
                release_state <= 3'h7;
              end else begin
                if(releaseDone) begin
                  release_state <= 3'h0;
                end else begin
                  if(s2_probe) begin
                    if(T_4375) begin
                      release_state <= 3'h5;
                    end else begin
                      if(T_4370) begin
                        release_state <= 3'h4;
                      end else begin
                        if(T_4196) begin
                          release_state <= 3'h3;
                        end else begin
                          if(T_4356) begin
                            release_state <= 3'h2;
                          end
                        end
                      end
                    end
                  end else begin
                    if(T_4356) begin
                      release_state <= 3'h2;
                    end
                  end
                end
              end
            end else begin
              if(releaseDone) begin
                release_state <= 3'h0;
              end else begin
                if(s2_probe) begin
                  if(T_4375) begin
                    release_state <= 3'h5;
                  end else begin
                    if(T_4370) begin
                      release_state <= 3'h4;
                    end else begin
                      if(T_4196) begin
                        release_state <= 3'h3;
                      end else begin
                        if(T_4356) begin
                          release_state <= 3'h2;
                        end
                      end
                    end
                  end
                end else begin
                  if(T_4356) begin
                    release_state <= 3'h2;
                  end
                end
              end
            end
          end
        end else begin
          if(T_4383) begin
            if(releaseDone) begin
              release_state <= 3'h7;
            end else begin
              if(releaseDone) begin
                release_state <= 3'h0;
              end else begin
                if(s2_probe) begin
                  if(T_4375) begin
                    release_state <= 3'h5;
                  end else begin
                    if(T_4370) begin
                      release_state <= 3'h4;
                    end else begin
                      if(T_4196) begin
                        release_state <= 3'h3;
                      end else begin
                        release_state <= GEN_79;
                      end
                    end
                  end
                end else begin
                  release_state <= GEN_79;
                end
              end
            end
          end else begin
            if(releaseDone) begin
              release_state <= 3'h0;
            end else begin
              if(s2_probe) begin
                if(T_4375) begin
                  release_state <= 3'h5;
                end else begin
                  if(T_4370) begin
                    release_state <= 3'h4;
                  end else begin
                    if(T_4196) begin
                      release_state <= 3'h3;
                    end else begin
                      release_state <= GEN_79;
                    end
                  end
                end
              end else begin
                release_state <= GEN_79;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      pstore2_valid <= T_2989;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    if(reset) begin
      s2_probe <= 1'h0;
    end else begin
      s2_probe <= s1_probe;
    end
    if(1'h0) begin
    end else begin
      T_2591 <= T_2257;
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        s2_req_addr <= {{8'd0}, s1_paddr};
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        s2_req_tag <= s1_req_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        s2_req_cmd <= s1_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        s2_req_typ <= s1_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        s2_req_phys <= s1_req_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        s2_req_data <= s1_req_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        s2_uncached <= T_2661;
      end
    end
    if(1'h0) begin
    end else begin
      s2_flush_valid <= s1_flush_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_mem_grant_valid) begin
        if(grantIsUncached) begin
          s2_data <= io_mem_grant_bits_data;
        end else begin
          if(T_2678) begin
            s2_data <= data_io_resp_0;
          end
        end
      end else begin
        if(T_2678) begin
          s2_data <= data_io_resp_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_probe) begin
        s2_probe_way <= s1_hit_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_probe) begin
        s2_probe_state_state <= s1_hit_state_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_valid_not_nacked) begin
        s2_hit_way <= s1_hit_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_valid_not_nacked) begin
        s2_hit_state_state <= s1_hit_state_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        T_2756 <= s1_victim_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        s2_victim_tag <= GEN_0_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        T_2766_state <= GEN_1_coh_state;
      end
    end
    if(reset) begin
      lrscCount <= 5'h0;
    end else begin
      if(T_2907) begin
        lrscCount <= 5'h0;
      end else begin
        if(lrscValid) begin
          lrscCount <= T_2905;
        end else begin
          if(T_2900) begin
            lrscCount <= 5'h1f;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2900) begin
        lrscAddr <= T_2895;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2909) begin
        pstore1_cmd <= s1_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2909) begin
        pstore1_typ <= s1_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2909) begin
        pstore1_addr <= s1_paddr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2909) begin
        pstore1_data <= io_cpu_s1_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2909) begin
        pstore1_way <= s1_hit_way;
      end
    end
    if(1'h0) begin
    end else begin
      T_2970 <= T_2983;
    end
    if(1'h0) begin
    end else begin
      if(advance_pstore1) begin
        pstore2_addr <= pstore1_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(advance_pstore1) begin
        pstore2_way <= pstore1_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(advance_pstore1) begin
        pstore2_storegen_data <= pstore1_storegen_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(advance_pstore1) begin
        pstore2_storegen_mask <= T_3029;
      end
    end
    if(reset) begin
      refillCount <= 3'h0;
    end else begin
      if(T_3743) begin
        refillCount <= T_3749;
      end
    end
    if(reset) begin
      writebackCount <= 3'h0;
    end else begin
      if(T_3911) begin
        writebackCount <= T_3917;
      end
    end
    if(1'h0) begin
    end else begin
      s1_release_data_valid <= T_3924;
    end
    if(1'h0) begin
    end else begin
      s2_release_data_valid <= T_3927;
    end
    if(1'h0) begin
    end else begin
      doUncachedResp <= io_cpu_replay_next;
    end
    if(reset) begin
      flushed <= 1'h1;
    end else begin
      if(flushing) begin
        if(s2_flush_valid) begin
          if(T_4547) begin
            flushed <= 1'h1;
          end else begin
            if(T_4521) begin
              flushed <= 1'h0;
            end
          end
        end else begin
          if(T_4521) begin
            flushed <= 1'h0;
          end
        end
      end else begin
        if(T_4521) begin
          flushed <= 1'h0;
        end
      end
    end
    if(reset) begin
      flushing <= 1'h0;
    end else begin
      if(flushing) begin
        if(T_4556) begin
          flushing <= 1'h0;
        end else begin
          if(T_4524) begin
            if(T_4526) begin
              flushing <= T_2748;
            end
          end
        end
      end else begin
        if(T_4524) begin
          if(T_4526) begin
            flushing <= T_2748;
          end
        end
      end
    end
    if(reset) begin
      T_4517 <= 6'h0;
    end else begin
      if(flushing) begin
        if(s2_flush_valid) begin
          T_4517 <= T_4550;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2978) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:214 assert(!s2_store_valid || !pstore1_held)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_2978) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_uncached & T_3715) begin
          $fwrite(32'h80000002,"Assertion failed: cache hit on uncached access\n    at dcache.scala:277 assert(!s2_valid_masked || !s2_hit_state.isValid(), \"cache hit on uncached access\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (s2_uncached & T_3715) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_mem_grant_valid & T_3740) begin
          $fwrite(32'h80000002,"Assertion failed: unexpected grant\n    at dcache.scala:293 assert(grant_wait || grantIsVoluntary && release_ack_wait, \"unexpected grant\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_mem_grant_valid & T_3740) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_3760) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:304 assert(dataArb.io.in(1).ready || !dataArb.io.in(1).valid)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_3760) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_3772) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:312 assert(!metaWriteArb.io.in(1).valid || metaWriteArb.io.in(1).ready)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_3772) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fq_io_enq_valid & T_3891) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:322 when (fq.io.enq.valid) { assert(fq.io.enq.ready) }\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (fq_io_enq_valid & T_3891) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_4356 & T_4363) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:348 assert(!(s2_valid && s2_hit_state.isValid()))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_4356 & T_4363) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doUncachedResp & T_4424) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:405 assert(!s2_valid_hit)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doUncachedResp & T_4424) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOArbiter(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input   io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output  io_in_0_grant_bits_client_xact_id,
  output [1:0] io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output  io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [10:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input   io_out_grant_bits_client_xact_id,
  input  [1:0] io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module HellaCacheArbiter(
  input   clk,
  input   reset,
  output  io_requestor_0_req_ready,
  input   io_requestor_0_req_valid,
  input  [39:0] io_requestor_0_req_bits_addr,
  input  [5:0] io_requestor_0_req_bits_tag,
  input  [4:0] io_requestor_0_req_bits_cmd,
  input  [2:0] io_requestor_0_req_bits_typ,
  input   io_requestor_0_req_bits_phys,
  input  [63:0] io_requestor_0_req_bits_data,
  input   io_requestor_0_s1_kill,
  input  [63:0] io_requestor_0_s1_data,
  output  io_requestor_0_s2_nack,
  output  io_requestor_0_resp_valid,
  output [39:0] io_requestor_0_resp_bits_addr,
  output [5:0] io_requestor_0_resp_bits_tag,
  output [4:0] io_requestor_0_resp_bits_cmd,
  output [2:0] io_requestor_0_resp_bits_typ,
  output [63:0] io_requestor_0_resp_bits_data,
  output  io_requestor_0_resp_bits_replay,
  output  io_requestor_0_resp_bits_has_data,
  output [63:0] io_requestor_0_resp_bits_data_word_bypass,
  output [63:0] io_requestor_0_resp_bits_store_data,
  output  io_requestor_0_replay_next,
  output  io_requestor_0_xcpt_ma_ld,
  output  io_requestor_0_xcpt_ma_st,
  output  io_requestor_0_xcpt_pf_ld,
  output  io_requestor_0_xcpt_pf_st,
  input   io_requestor_0_invalidate_lr,
  output  io_requestor_0_ordered,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [5:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [2:0] io_mem_req_bits_typ,
  output  io_mem_req_bits_phys,
  output [63:0] io_mem_req_bits_data,
  output  io_mem_s1_kill,
  output [63:0] io_mem_s1_data,
  input   io_mem_s2_nack,
  input   io_mem_resp_valid,
  input  [39:0] io_mem_resp_bits_addr,
  input  [5:0] io_mem_resp_bits_tag,
  input  [4:0] io_mem_resp_bits_cmd,
  input  [2:0] io_mem_resp_bits_typ,
  input  [63:0] io_mem_resp_bits_data,
  input   io_mem_resp_bits_replay,
  input   io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input  [63:0] io_mem_resp_bits_store_data,
  input   io_mem_replay_next,
  input   io_mem_xcpt_ma_ld,
  input   io_mem_xcpt_ma_st,
  input   io_mem_xcpt_pf_ld,
  input   io_mem_xcpt_pf_st,
  output  io_mem_invalidate_lr,
  input   io_mem_ordered
);
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_0_s2_nack = io_mem_s2_nack;
  assign io_requestor_0_resp_valid = io_mem_resp_valid;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_tag = io_mem_resp_bits_tag;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_replay = io_mem_resp_bits_replay;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_replay_next = io_mem_replay_next;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_mem_req_valid = io_requestor_0_req_valid;
  assign io_mem_req_bits_addr = io_requestor_0_req_bits_addr;
  assign io_mem_req_bits_tag = io_requestor_0_req_bits_tag;
  assign io_mem_req_bits_cmd = io_requestor_0_req_bits_cmd;
  assign io_mem_req_bits_typ = io_requestor_0_req_bits_typ;
  assign io_mem_req_bits_phys = io_requestor_0_req_bits_phys;
  assign io_mem_req_bits_data = io_requestor_0_req_bits_data;
  assign io_mem_s1_kill = io_requestor_0_s1_kill;
  assign io_mem_s1_data = io_requestor_0_s1_data;
  assign io_mem_invalidate_lr = io_requestor_0_invalidate_lr;
endmodule
module RocketTile(
  input   clk,
  input   reset,
  input   io_cached_0_acquire_ready,
  output  io_cached_0_acquire_valid,
  output [25:0] io_cached_0_acquire_bits_addr_block,
  output  io_cached_0_acquire_bits_client_xact_id,
  output [2:0] io_cached_0_acquire_bits_addr_beat,
  output  io_cached_0_acquire_bits_is_builtin_type,
  output [2:0] io_cached_0_acquire_bits_a_type,
  output [10:0] io_cached_0_acquire_bits_union,
  output [63:0] io_cached_0_acquire_bits_data,
  output  io_cached_0_probe_ready,
  input   io_cached_0_probe_valid,
  input  [25:0] io_cached_0_probe_bits_addr_block,
  input  [1:0] io_cached_0_probe_bits_p_type,
  input   io_cached_0_release_ready,
  output  io_cached_0_release_valid,
  output [2:0] io_cached_0_release_bits_addr_beat,
  output [25:0] io_cached_0_release_bits_addr_block,
  output  io_cached_0_release_bits_client_xact_id,
  output  io_cached_0_release_bits_voluntary,
  output [2:0] io_cached_0_release_bits_r_type,
  output [63:0] io_cached_0_release_bits_data,
  output  io_cached_0_grant_ready,
  input   io_cached_0_grant_valid,
  input  [2:0] io_cached_0_grant_bits_addr_beat,
  input   io_cached_0_grant_bits_client_xact_id,
  input  [1:0] io_cached_0_grant_bits_manager_xact_id,
  input   io_cached_0_grant_bits_is_builtin_type,
  input  [3:0] io_cached_0_grant_bits_g_type,
  input  [63:0] io_cached_0_grant_bits_data,
  input   io_cached_0_grant_bits_manager_id,
  input   io_cached_0_finish_ready,
  output  io_cached_0_finish_valid,
  output [1:0] io_cached_0_finish_bits_manager_xact_id,
  output  io_cached_0_finish_bits_manager_id,
  input   io_uncached_0_acquire_ready,
  output  io_uncached_0_acquire_valid,
  output [25:0] io_uncached_0_acquire_bits_addr_block,
  output  io_uncached_0_acquire_bits_client_xact_id,
  output [2:0] io_uncached_0_acquire_bits_addr_beat,
  output  io_uncached_0_acquire_bits_is_builtin_type,
  output [2:0] io_uncached_0_acquire_bits_a_type,
  output [10:0] io_uncached_0_acquire_bits_union,
  output [63:0] io_uncached_0_acquire_bits_data,
  output  io_uncached_0_grant_ready,
  input   io_uncached_0_grant_valid,
  input  [2:0] io_uncached_0_grant_bits_addr_beat,
  input   io_uncached_0_grant_bits_client_xact_id,
  input  [1:0] io_uncached_0_grant_bits_manager_xact_id,
  input   io_uncached_0_grant_bits_is_builtin_type,
  input  [3:0] io_uncached_0_grant_bits_g_type,
  input  [63:0] io_uncached_0_grant_bits_data,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip
);
  wire  core_clk;
  wire  core_reset;
  wire  core_io_prci_reset;
  wire  core_io_prci_id;
  wire  core_io_prci_interrupts_meip;
  wire  core_io_prci_interrupts_seip;
  wire  core_io_prci_interrupts_debug;
  wire  core_io_prci_interrupts_mtip;
  wire  core_io_prci_interrupts_msip;
  wire  core_io_imem_req_valid;
  wire [39:0] core_io_imem_req_bits_pc;
  wire  core_io_imem_req_bits_speculative;
  wire  core_io_imem_resp_ready;
  wire  core_io_imem_resp_valid;
  wire  core_io_imem_resp_bits_btb_valid;
  wire  core_io_imem_resp_bits_btb_bits_taken;
  wire [1:0] core_io_imem_resp_bits_btb_bits_mask;
  wire  core_io_imem_resp_bits_btb_bits_bridx;
  wire [38:0] core_io_imem_resp_bits_btb_bits_target;
  wire  core_io_imem_resp_bits_btb_bits_entry;
  wire  core_io_imem_resp_bits_btb_bits_bht_history;
  wire [1:0] core_io_imem_resp_bits_btb_bits_bht_value;
  wire [39:0] core_io_imem_resp_bits_pc;
  wire [31:0] core_io_imem_resp_bits_data;
  wire [1:0] core_io_imem_resp_bits_mask;
  wire  core_io_imem_resp_bits_xcpt_if;
  wire  core_io_imem_resp_bits_replay;
  wire  core_io_imem_btb_update_valid;
  wire  core_io_imem_btb_update_bits_prediction_valid;
  wire  core_io_imem_btb_update_bits_prediction_bits_taken;
  wire [1:0] core_io_imem_btb_update_bits_prediction_bits_mask;
  wire  core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire  core_io_imem_btb_update_bits_prediction_bits_entry;
  wire  core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] core_io_imem_btb_update_bits_pc;
  wire [38:0] core_io_imem_btb_update_bits_target;
  wire  core_io_imem_btb_update_bits_taken;
  wire  core_io_imem_btb_update_bits_isValid;
  wire  core_io_imem_btb_update_bits_isJump;
  wire  core_io_imem_btb_update_bits_isReturn;
  wire [38:0] core_io_imem_btb_update_bits_br_pc;
  wire  core_io_imem_bht_update_valid;
  wire  core_io_imem_bht_update_bits_prediction_valid;
  wire  core_io_imem_bht_update_bits_prediction_bits_taken;
  wire [1:0] core_io_imem_bht_update_bits_prediction_bits_mask;
  wire  core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire  core_io_imem_bht_update_bits_prediction_bits_entry;
  wire  core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] core_io_imem_bht_update_bits_pc;
  wire  core_io_imem_bht_update_bits_taken;
  wire  core_io_imem_bht_update_bits_mispredict;
  wire  core_io_imem_ras_update_valid;
  wire  core_io_imem_ras_update_bits_isCall;
  wire  core_io_imem_ras_update_bits_isReturn;
  wire [38:0] core_io_imem_ras_update_bits_returnAddr;
  wire  core_io_imem_ras_update_bits_prediction_valid;
  wire  core_io_imem_ras_update_bits_prediction_bits_taken;
  wire [1:0] core_io_imem_ras_update_bits_prediction_bits_mask;
  wire  core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire  core_io_imem_ras_update_bits_prediction_bits_entry;
  wire  core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire  core_io_imem_flush_icache;
  wire  core_io_imem_flush_tlb;
  wire [39:0] core_io_imem_npc;
  wire  core_io_dmem_req_ready;
  wire  core_io_dmem_req_valid;
  wire [39:0] core_io_dmem_req_bits_addr;
  wire [5:0] core_io_dmem_req_bits_tag;
  wire [4:0] core_io_dmem_req_bits_cmd;
  wire [2:0] core_io_dmem_req_bits_typ;
  wire  core_io_dmem_req_bits_phys;
  wire [63:0] core_io_dmem_req_bits_data;
  wire  core_io_dmem_s1_kill;
  wire [63:0] core_io_dmem_s1_data;
  wire  core_io_dmem_s2_nack;
  wire  core_io_dmem_resp_valid;
  wire [39:0] core_io_dmem_resp_bits_addr;
  wire [5:0] core_io_dmem_resp_bits_tag;
  wire [4:0] core_io_dmem_resp_bits_cmd;
  wire [2:0] core_io_dmem_resp_bits_typ;
  wire [63:0] core_io_dmem_resp_bits_data;
  wire  core_io_dmem_resp_bits_replay;
  wire  core_io_dmem_resp_bits_has_data;
  wire [63:0] core_io_dmem_resp_bits_data_word_bypass;
  wire [63:0] core_io_dmem_resp_bits_store_data;
  wire  core_io_dmem_replay_next;
  wire  core_io_dmem_xcpt_ma_ld;
  wire  core_io_dmem_xcpt_ma_st;
  wire  core_io_dmem_xcpt_pf_ld;
  wire  core_io_dmem_xcpt_pf_st;
  wire  core_io_dmem_invalidate_lr;
  wire  core_io_dmem_ordered;
  wire [6:0] core_io_ptw_ptbr_asid;
  wire [37:0] core_io_ptw_ptbr_ppn;
  wire  core_io_ptw_invalidate;
  wire  core_io_ptw_status_debug;
  wire [1:0] core_io_ptw_status_prv;
  wire  core_io_ptw_status_sd;
  wire [30:0] core_io_ptw_status_zero3;
  wire  core_io_ptw_status_sd_rv32;
  wire [1:0] core_io_ptw_status_zero2;
  wire [4:0] core_io_ptw_status_vm;
  wire [3:0] core_io_ptw_status_zero1;
  wire  core_io_ptw_status_mxr;
  wire  core_io_ptw_status_pum;
  wire  core_io_ptw_status_mprv;
  wire [1:0] core_io_ptw_status_xs;
  wire [1:0] core_io_ptw_status_fs;
  wire [1:0] core_io_ptw_status_mpp;
  wire [1:0] core_io_ptw_status_hpp;
  wire  core_io_ptw_status_spp;
  wire  core_io_ptw_status_mpie;
  wire  core_io_ptw_status_hpie;
  wire  core_io_ptw_status_spie;
  wire  core_io_ptw_status_upie;
  wire  core_io_ptw_status_mie;
  wire  core_io_ptw_status_hie;
  wire  core_io_ptw_status_sie;
  wire  core_io_ptw_status_uie;
  wire [31:0] core_io_fpu_inst;
  wire [63:0] core_io_fpu_fromint_data;
  wire [2:0] core_io_fpu_fcsr_rm;
  wire  core_io_fpu_fcsr_flags_valid;
  wire [4:0] core_io_fpu_fcsr_flags_bits;
  wire [63:0] core_io_fpu_store_data;
  wire [63:0] core_io_fpu_toint_data;
  wire  core_io_fpu_dmem_resp_val;
  wire [2:0] core_io_fpu_dmem_resp_type;
  wire [4:0] core_io_fpu_dmem_resp_tag;
  wire [63:0] core_io_fpu_dmem_resp_data;
  wire  core_io_fpu_valid;
  wire  core_io_fpu_fcsr_rdy;
  wire  core_io_fpu_nack_mem;
  wire  core_io_fpu_illegal_rm;
  wire  core_io_fpu_killx;
  wire  core_io_fpu_killm;
  wire [4:0] core_io_fpu_dec_cmd;
  wire  core_io_fpu_dec_ldst;
  wire  core_io_fpu_dec_wen;
  wire  core_io_fpu_dec_ren1;
  wire  core_io_fpu_dec_ren2;
  wire  core_io_fpu_dec_ren3;
  wire  core_io_fpu_dec_swap12;
  wire  core_io_fpu_dec_swap23;
  wire  core_io_fpu_dec_single;
  wire  core_io_fpu_dec_fromint;
  wire  core_io_fpu_dec_toint;
  wire  core_io_fpu_dec_fastpipe;
  wire  core_io_fpu_dec_fma;
  wire  core_io_fpu_dec_div;
  wire  core_io_fpu_dec_sqrt;
  wire  core_io_fpu_dec_round;
  wire  core_io_fpu_dec_wflags;
  wire  core_io_fpu_sboard_set;
  wire  core_io_fpu_sboard_clr;
  wire [4:0] core_io_fpu_sboard_clra;
  wire  core_io_fpu_cp_req_ready;
  wire  core_io_fpu_cp_req_valid;
  wire [4:0] core_io_fpu_cp_req_bits_cmd;
  wire  core_io_fpu_cp_req_bits_ldst;
  wire  core_io_fpu_cp_req_bits_wen;
  wire  core_io_fpu_cp_req_bits_ren1;
  wire  core_io_fpu_cp_req_bits_ren2;
  wire  core_io_fpu_cp_req_bits_ren3;
  wire  core_io_fpu_cp_req_bits_swap12;
  wire  core_io_fpu_cp_req_bits_swap23;
  wire  core_io_fpu_cp_req_bits_single;
  wire  core_io_fpu_cp_req_bits_fromint;
  wire  core_io_fpu_cp_req_bits_toint;
  wire  core_io_fpu_cp_req_bits_fastpipe;
  wire  core_io_fpu_cp_req_bits_fma;
  wire  core_io_fpu_cp_req_bits_div;
  wire  core_io_fpu_cp_req_bits_sqrt;
  wire  core_io_fpu_cp_req_bits_round;
  wire  core_io_fpu_cp_req_bits_wflags;
  wire [2:0] core_io_fpu_cp_req_bits_rm;
  wire [1:0] core_io_fpu_cp_req_bits_typ;
  wire [64:0] core_io_fpu_cp_req_bits_in1;
  wire [64:0] core_io_fpu_cp_req_bits_in2;
  wire [64:0] core_io_fpu_cp_req_bits_in3;
  wire  core_io_fpu_cp_resp_ready;
  wire  core_io_fpu_cp_resp_valid;
  wire [64:0] core_io_fpu_cp_resp_bits_data;
  wire [4:0] core_io_fpu_cp_resp_bits_exc;
  wire  core_io_rocc_cmd_ready;
  wire  core_io_rocc_cmd_valid;
  wire [6:0] core_io_rocc_cmd_bits_inst_funct;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs1;
  wire  core_io_rocc_cmd_bits_inst_xd;
  wire  core_io_rocc_cmd_bits_inst_xs1;
  wire  core_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rd;
  wire [6:0] core_io_rocc_cmd_bits_inst_opcode;
  wire [63:0] core_io_rocc_cmd_bits_rs1;
  wire [63:0] core_io_rocc_cmd_bits_rs2;
  wire  core_io_rocc_cmd_bits_status_debug;
  wire [1:0] core_io_rocc_cmd_bits_status_prv;
  wire  core_io_rocc_cmd_bits_status_sd;
  wire [30:0] core_io_rocc_cmd_bits_status_zero3;
  wire  core_io_rocc_cmd_bits_status_sd_rv32;
  wire [1:0] core_io_rocc_cmd_bits_status_zero2;
  wire [4:0] core_io_rocc_cmd_bits_status_vm;
  wire [3:0] core_io_rocc_cmd_bits_status_zero1;
  wire  core_io_rocc_cmd_bits_status_mxr;
  wire  core_io_rocc_cmd_bits_status_pum;
  wire  core_io_rocc_cmd_bits_status_mprv;
  wire [1:0] core_io_rocc_cmd_bits_status_xs;
  wire [1:0] core_io_rocc_cmd_bits_status_fs;
  wire [1:0] core_io_rocc_cmd_bits_status_mpp;
  wire [1:0] core_io_rocc_cmd_bits_status_hpp;
  wire  core_io_rocc_cmd_bits_status_spp;
  wire  core_io_rocc_cmd_bits_status_mpie;
  wire  core_io_rocc_cmd_bits_status_hpie;
  wire  core_io_rocc_cmd_bits_status_spie;
  wire  core_io_rocc_cmd_bits_status_upie;
  wire  core_io_rocc_cmd_bits_status_mie;
  wire  core_io_rocc_cmd_bits_status_hie;
  wire  core_io_rocc_cmd_bits_status_sie;
  wire  core_io_rocc_cmd_bits_status_uie;
  wire  core_io_rocc_resp_ready;
  wire  core_io_rocc_resp_valid;
  wire [4:0] core_io_rocc_resp_bits_rd;
  wire [63:0] core_io_rocc_resp_bits_data;
  wire  core_io_rocc_mem_req_ready;
  wire  core_io_rocc_mem_req_valid;
  wire [39:0] core_io_rocc_mem_req_bits_addr;
  wire [5:0] core_io_rocc_mem_req_bits_tag;
  wire [4:0] core_io_rocc_mem_req_bits_cmd;
  wire [2:0] core_io_rocc_mem_req_bits_typ;
  wire  core_io_rocc_mem_req_bits_phys;
  wire [63:0] core_io_rocc_mem_req_bits_data;
  wire  core_io_rocc_mem_s1_kill;
  wire [63:0] core_io_rocc_mem_s1_data;
  wire  core_io_rocc_mem_s2_nack;
  wire  core_io_rocc_mem_resp_valid;
  wire [39:0] core_io_rocc_mem_resp_bits_addr;
  wire [5:0] core_io_rocc_mem_resp_bits_tag;
  wire [4:0] core_io_rocc_mem_resp_bits_cmd;
  wire [2:0] core_io_rocc_mem_resp_bits_typ;
  wire [63:0] core_io_rocc_mem_resp_bits_data;
  wire  core_io_rocc_mem_resp_bits_replay;
  wire  core_io_rocc_mem_resp_bits_has_data;
  wire [63:0] core_io_rocc_mem_resp_bits_data_word_bypass;
  wire [63:0] core_io_rocc_mem_resp_bits_store_data;
  wire  core_io_rocc_mem_replay_next;
  wire  core_io_rocc_mem_xcpt_ma_ld;
  wire  core_io_rocc_mem_xcpt_ma_st;
  wire  core_io_rocc_mem_xcpt_pf_ld;
  wire  core_io_rocc_mem_xcpt_pf_st;
  wire  core_io_rocc_mem_invalidate_lr;
  wire  core_io_rocc_mem_ordered;
  wire  core_io_rocc_busy;
  wire  core_io_rocc_interrupt;
  wire  core_io_rocc_autl_acquire_ready;
  wire  core_io_rocc_autl_acquire_valid;
  wire [25:0] core_io_rocc_autl_acquire_bits_addr_block;
  wire  core_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] core_io_rocc_autl_acquire_bits_addr_beat;
  wire  core_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] core_io_rocc_autl_acquire_bits_a_type;
  wire [10:0] core_io_rocc_autl_acquire_bits_union;
  wire [63:0] core_io_rocc_autl_acquire_bits_data;
  wire  core_io_rocc_autl_grant_ready;
  wire  core_io_rocc_autl_grant_valid;
  wire [2:0] core_io_rocc_autl_grant_bits_addr_beat;
  wire  core_io_rocc_autl_grant_bits_client_xact_id;
  wire [1:0] core_io_rocc_autl_grant_bits_manager_xact_id;
  wire  core_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] core_io_rocc_autl_grant_bits_g_type;
  wire [63:0] core_io_rocc_autl_grant_bits_data;
  wire  core_io_rocc_fpu_req_ready;
  wire  core_io_rocc_fpu_req_valid;
  wire [4:0] core_io_rocc_fpu_req_bits_cmd;
  wire  core_io_rocc_fpu_req_bits_ldst;
  wire  core_io_rocc_fpu_req_bits_wen;
  wire  core_io_rocc_fpu_req_bits_ren1;
  wire  core_io_rocc_fpu_req_bits_ren2;
  wire  core_io_rocc_fpu_req_bits_ren3;
  wire  core_io_rocc_fpu_req_bits_swap12;
  wire  core_io_rocc_fpu_req_bits_swap23;
  wire  core_io_rocc_fpu_req_bits_single;
  wire  core_io_rocc_fpu_req_bits_fromint;
  wire  core_io_rocc_fpu_req_bits_toint;
  wire  core_io_rocc_fpu_req_bits_fastpipe;
  wire  core_io_rocc_fpu_req_bits_fma;
  wire  core_io_rocc_fpu_req_bits_div;
  wire  core_io_rocc_fpu_req_bits_sqrt;
  wire  core_io_rocc_fpu_req_bits_round;
  wire  core_io_rocc_fpu_req_bits_wflags;
  wire [2:0] core_io_rocc_fpu_req_bits_rm;
  wire [1:0] core_io_rocc_fpu_req_bits_typ;
  wire [64:0] core_io_rocc_fpu_req_bits_in1;
  wire [64:0] core_io_rocc_fpu_req_bits_in2;
  wire [64:0] core_io_rocc_fpu_req_bits_in3;
  wire  core_io_rocc_fpu_resp_ready;
  wire  core_io_rocc_fpu_resp_valid;
  wire [64:0] core_io_rocc_fpu_resp_bits_data;
  wire [4:0] core_io_rocc_fpu_resp_bits_exc;
  wire  core_io_rocc_exception;
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_cpu_req_valid;
  wire [39:0] icache_io_cpu_req_bits_pc;
  wire  icache_io_cpu_req_bits_speculative;
  wire  icache_io_cpu_resp_ready;
  wire  icache_io_cpu_resp_valid;
  wire  icache_io_cpu_resp_bits_btb_valid;
  wire  icache_io_cpu_resp_bits_btb_bits_taken;
  wire [1:0] icache_io_cpu_resp_bits_btb_bits_mask;
  wire  icache_io_cpu_resp_bits_btb_bits_bridx;
  wire [38:0] icache_io_cpu_resp_bits_btb_bits_target;
  wire  icache_io_cpu_resp_bits_btb_bits_entry;
  wire  icache_io_cpu_resp_bits_btb_bits_bht_history;
  wire [1:0] icache_io_cpu_resp_bits_btb_bits_bht_value;
  wire [39:0] icache_io_cpu_resp_bits_pc;
  wire [31:0] icache_io_cpu_resp_bits_data;
  wire [1:0] icache_io_cpu_resp_bits_mask;
  wire  icache_io_cpu_resp_bits_xcpt_if;
  wire  icache_io_cpu_resp_bits_replay;
  wire  icache_io_cpu_btb_update_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_taken;
  wire [1:0] icache_io_cpu_btb_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_btb_update_bits_prediction_bits_target;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_entry;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] icache_io_cpu_btb_update_bits_pc;
  wire [38:0] icache_io_cpu_btb_update_bits_target;
  wire  icache_io_cpu_btb_update_bits_taken;
  wire  icache_io_cpu_btb_update_bits_isValid;
  wire  icache_io_cpu_btb_update_bits_isJump;
  wire  icache_io_cpu_btb_update_bits_isReturn;
  wire [38:0] icache_io_cpu_btb_update_bits_br_pc;
  wire  icache_io_cpu_bht_update_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_taken;
  wire [1:0] icache_io_cpu_bht_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_bht_update_bits_prediction_bits_target;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_entry;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] icache_io_cpu_bht_update_bits_pc;
  wire  icache_io_cpu_bht_update_bits_taken;
  wire  icache_io_cpu_bht_update_bits_mispredict;
  wire  icache_io_cpu_ras_update_valid;
  wire  icache_io_cpu_ras_update_bits_isCall;
  wire  icache_io_cpu_ras_update_bits_isReturn;
  wire [38:0] icache_io_cpu_ras_update_bits_returnAddr;
  wire  icache_io_cpu_ras_update_bits_prediction_valid;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_taken;
  wire [1:0] icache_io_cpu_ras_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_ras_update_bits_prediction_bits_target;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_entry;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_ras_update_bits_prediction_bits_bht_value;
  wire  icache_io_cpu_flush_icache;
  wire  icache_io_cpu_flush_tlb;
  wire [39:0] icache_io_cpu_npc;
  wire  icache_io_ptw_req_ready;
  wire  icache_io_ptw_req_valid;
  wire [1:0] icache_io_ptw_req_bits_prv;
  wire  icache_io_ptw_req_bits_pum;
  wire  icache_io_ptw_req_bits_mxr;
  wire [26:0] icache_io_ptw_req_bits_addr;
  wire  icache_io_ptw_req_bits_store;
  wire  icache_io_ptw_req_bits_fetch;
  wire  icache_io_ptw_resp_valid;
  wire [15:0] icache_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] icache_io_ptw_resp_bits_pte_ppn;
  wire [1:0] icache_io_ptw_resp_bits_pte_reserved_for_software;
  wire  icache_io_ptw_resp_bits_pte_d;
  wire  icache_io_ptw_resp_bits_pte_a;
  wire  icache_io_ptw_resp_bits_pte_g;
  wire  icache_io_ptw_resp_bits_pte_u;
  wire  icache_io_ptw_resp_bits_pte_x;
  wire  icache_io_ptw_resp_bits_pte_w;
  wire  icache_io_ptw_resp_bits_pte_r;
  wire  icache_io_ptw_resp_bits_pte_v;
  wire [6:0] icache_io_ptw_ptbr_asid;
  wire [37:0] icache_io_ptw_ptbr_ppn;
  wire  icache_io_ptw_invalidate;
  wire  icache_io_ptw_status_debug;
  wire [1:0] icache_io_ptw_status_prv;
  wire  icache_io_ptw_status_sd;
  wire [30:0] icache_io_ptw_status_zero3;
  wire  icache_io_ptw_status_sd_rv32;
  wire [1:0] icache_io_ptw_status_zero2;
  wire [4:0] icache_io_ptw_status_vm;
  wire [3:0] icache_io_ptw_status_zero1;
  wire  icache_io_ptw_status_mxr;
  wire  icache_io_ptw_status_pum;
  wire  icache_io_ptw_status_mprv;
  wire [1:0] icache_io_ptw_status_xs;
  wire [1:0] icache_io_ptw_status_fs;
  wire [1:0] icache_io_ptw_status_mpp;
  wire [1:0] icache_io_ptw_status_hpp;
  wire  icache_io_ptw_status_spp;
  wire  icache_io_ptw_status_mpie;
  wire  icache_io_ptw_status_hpie;
  wire  icache_io_ptw_status_spie;
  wire  icache_io_ptw_status_upie;
  wire  icache_io_ptw_status_mie;
  wire  icache_io_ptw_status_hie;
  wire  icache_io_ptw_status_sie;
  wire  icache_io_ptw_status_uie;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire  icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [10:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire  icache_io_mem_grant_bits_client_xact_id;
  wire [1:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  DCache_1_clk;
  wire  DCache_1_reset;
  wire  DCache_1_io_cpu_req_ready;
  wire  DCache_1_io_cpu_req_valid;
  wire [39:0] DCache_1_io_cpu_req_bits_addr;
  wire [5:0] DCache_1_io_cpu_req_bits_tag;
  wire [4:0] DCache_1_io_cpu_req_bits_cmd;
  wire [2:0] DCache_1_io_cpu_req_bits_typ;
  wire  DCache_1_io_cpu_req_bits_phys;
  wire [63:0] DCache_1_io_cpu_req_bits_data;
  wire  DCache_1_io_cpu_s1_kill;
  wire [63:0] DCache_1_io_cpu_s1_data;
  wire  DCache_1_io_cpu_s2_nack;
  wire  DCache_1_io_cpu_resp_valid;
  wire [39:0] DCache_1_io_cpu_resp_bits_addr;
  wire [5:0] DCache_1_io_cpu_resp_bits_tag;
  wire [4:0] DCache_1_io_cpu_resp_bits_cmd;
  wire [2:0] DCache_1_io_cpu_resp_bits_typ;
  wire [63:0] DCache_1_io_cpu_resp_bits_data;
  wire  DCache_1_io_cpu_resp_bits_replay;
  wire  DCache_1_io_cpu_resp_bits_has_data;
  wire [63:0] DCache_1_io_cpu_resp_bits_data_word_bypass;
  wire [63:0] DCache_1_io_cpu_resp_bits_store_data;
  wire  DCache_1_io_cpu_replay_next;
  wire  DCache_1_io_cpu_xcpt_ma_ld;
  wire  DCache_1_io_cpu_xcpt_ma_st;
  wire  DCache_1_io_cpu_xcpt_pf_ld;
  wire  DCache_1_io_cpu_xcpt_pf_st;
  wire  DCache_1_io_cpu_invalidate_lr;
  wire  DCache_1_io_cpu_ordered;
  wire  DCache_1_io_ptw_req_ready;
  wire  DCache_1_io_ptw_req_valid;
  wire [1:0] DCache_1_io_ptw_req_bits_prv;
  wire  DCache_1_io_ptw_req_bits_pum;
  wire  DCache_1_io_ptw_req_bits_mxr;
  wire [26:0] DCache_1_io_ptw_req_bits_addr;
  wire  DCache_1_io_ptw_req_bits_store;
  wire  DCache_1_io_ptw_req_bits_fetch;
  wire  DCache_1_io_ptw_resp_valid;
  wire [15:0] DCache_1_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] DCache_1_io_ptw_resp_bits_pte_ppn;
  wire [1:0] DCache_1_io_ptw_resp_bits_pte_reserved_for_software;
  wire  DCache_1_io_ptw_resp_bits_pte_d;
  wire  DCache_1_io_ptw_resp_bits_pte_a;
  wire  DCache_1_io_ptw_resp_bits_pte_g;
  wire  DCache_1_io_ptw_resp_bits_pte_u;
  wire  DCache_1_io_ptw_resp_bits_pte_x;
  wire  DCache_1_io_ptw_resp_bits_pte_w;
  wire  DCache_1_io_ptw_resp_bits_pte_r;
  wire  DCache_1_io_ptw_resp_bits_pte_v;
  wire [6:0] DCache_1_io_ptw_ptbr_asid;
  wire [37:0] DCache_1_io_ptw_ptbr_ppn;
  wire  DCache_1_io_ptw_invalidate;
  wire  DCache_1_io_ptw_status_debug;
  wire [1:0] DCache_1_io_ptw_status_prv;
  wire  DCache_1_io_ptw_status_sd;
  wire [30:0] DCache_1_io_ptw_status_zero3;
  wire  DCache_1_io_ptw_status_sd_rv32;
  wire [1:0] DCache_1_io_ptw_status_zero2;
  wire [4:0] DCache_1_io_ptw_status_vm;
  wire [3:0] DCache_1_io_ptw_status_zero1;
  wire  DCache_1_io_ptw_status_mxr;
  wire  DCache_1_io_ptw_status_pum;
  wire  DCache_1_io_ptw_status_mprv;
  wire [1:0] DCache_1_io_ptw_status_xs;
  wire [1:0] DCache_1_io_ptw_status_fs;
  wire [1:0] DCache_1_io_ptw_status_mpp;
  wire [1:0] DCache_1_io_ptw_status_hpp;
  wire  DCache_1_io_ptw_status_spp;
  wire  DCache_1_io_ptw_status_mpie;
  wire  DCache_1_io_ptw_status_hpie;
  wire  DCache_1_io_ptw_status_spie;
  wire  DCache_1_io_ptw_status_upie;
  wire  DCache_1_io_ptw_status_mie;
  wire  DCache_1_io_ptw_status_hie;
  wire  DCache_1_io_ptw_status_sie;
  wire  DCache_1_io_ptw_status_uie;
  wire  DCache_1_io_mem_acquire_ready;
  wire  DCache_1_io_mem_acquire_valid;
  wire [25:0] DCache_1_io_mem_acquire_bits_addr_block;
  wire  DCache_1_io_mem_acquire_bits_client_xact_id;
  wire [2:0] DCache_1_io_mem_acquire_bits_addr_beat;
  wire  DCache_1_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] DCache_1_io_mem_acquire_bits_a_type;
  wire [10:0] DCache_1_io_mem_acquire_bits_union;
  wire [63:0] DCache_1_io_mem_acquire_bits_data;
  wire  DCache_1_io_mem_probe_ready;
  wire  DCache_1_io_mem_probe_valid;
  wire [25:0] DCache_1_io_mem_probe_bits_addr_block;
  wire [1:0] DCache_1_io_mem_probe_bits_p_type;
  wire  DCache_1_io_mem_release_ready;
  wire  DCache_1_io_mem_release_valid;
  wire [2:0] DCache_1_io_mem_release_bits_addr_beat;
  wire [25:0] DCache_1_io_mem_release_bits_addr_block;
  wire  DCache_1_io_mem_release_bits_client_xact_id;
  wire  DCache_1_io_mem_release_bits_voluntary;
  wire [2:0] DCache_1_io_mem_release_bits_r_type;
  wire [63:0] DCache_1_io_mem_release_bits_data;
  wire  DCache_1_io_mem_grant_ready;
  wire  DCache_1_io_mem_grant_valid;
  wire [2:0] DCache_1_io_mem_grant_bits_addr_beat;
  wire  DCache_1_io_mem_grant_bits_client_xact_id;
  wire [1:0] DCache_1_io_mem_grant_bits_manager_xact_id;
  wire  DCache_1_io_mem_grant_bits_is_builtin_type;
  wire [3:0] DCache_1_io_mem_grant_bits_g_type;
  wire [63:0] DCache_1_io_mem_grant_bits_data;
  wire  DCache_1_io_mem_grant_bits_manager_id;
  wire  DCache_1_io_mem_finish_ready;
  wire  DCache_1_io_mem_finish_valid;
  wire [1:0] DCache_1_io_mem_finish_bits_manager_xact_id;
  wire  DCache_1_io_mem_finish_bits_manager_id;
  wire  uncachedArb_clk;
  wire  uncachedArb_reset;
  wire  uncachedArb_io_in_0_acquire_ready;
  wire  uncachedArb_io_in_0_acquire_valid;
  wire [25:0] uncachedArb_io_in_0_acquire_bits_addr_block;
  wire  uncachedArb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_addr_beat;
  wire  uncachedArb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_a_type;
  wire [10:0] uncachedArb_io_in_0_acquire_bits_union;
  wire [63:0] uncachedArb_io_in_0_acquire_bits_data;
  wire  uncachedArb_io_in_0_grant_ready;
  wire  uncachedArb_io_in_0_grant_valid;
  wire [2:0] uncachedArb_io_in_0_grant_bits_addr_beat;
  wire  uncachedArb_io_in_0_grant_bits_client_xact_id;
  wire [1:0] uncachedArb_io_in_0_grant_bits_manager_xact_id;
  wire  uncachedArb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_in_0_grant_bits_g_type;
  wire [63:0] uncachedArb_io_in_0_grant_bits_data;
  wire  uncachedArb_io_out_acquire_ready;
  wire  uncachedArb_io_out_acquire_valid;
  wire [25:0] uncachedArb_io_out_acquire_bits_addr_block;
  wire  uncachedArb_io_out_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_out_acquire_bits_addr_beat;
  wire  uncachedArb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_out_acquire_bits_a_type;
  wire [10:0] uncachedArb_io_out_acquire_bits_union;
  wire [63:0] uncachedArb_io_out_acquire_bits_data;
  wire  uncachedArb_io_out_grant_ready;
  wire  uncachedArb_io_out_grant_valid;
  wire [2:0] uncachedArb_io_out_grant_bits_addr_beat;
  wire  uncachedArb_io_out_grant_bits_client_xact_id;
  wire [1:0] uncachedArb_io_out_grant_bits_manager_xact_id;
  wire  uncachedArb_io_out_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_out_grant_bits_g_type;
  wire [63:0] uncachedArb_io_out_grant_bits_data;
  wire  dcArb_clk;
  wire  dcArb_reset;
  wire  dcArb_io_requestor_0_req_ready;
  wire  dcArb_io_requestor_0_req_valid;
  wire [39:0] dcArb_io_requestor_0_req_bits_addr;
  wire [5:0] dcArb_io_requestor_0_req_bits_tag;
  wire [4:0] dcArb_io_requestor_0_req_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_req_bits_typ;
  wire  dcArb_io_requestor_0_req_bits_phys;
  wire [63:0] dcArb_io_requestor_0_req_bits_data;
  wire  dcArb_io_requestor_0_s1_kill;
  wire [63:0] dcArb_io_requestor_0_s1_data;
  wire  dcArb_io_requestor_0_s2_nack;
  wire  dcArb_io_requestor_0_resp_valid;
  wire [39:0] dcArb_io_requestor_0_resp_bits_addr;
  wire [5:0] dcArb_io_requestor_0_resp_bits_tag;
  wire [4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire [63:0] dcArb_io_requestor_0_resp_bits_data;
  wire  dcArb_io_requestor_0_resp_bits_replay;
  wire  dcArb_io_requestor_0_resp_bits_has_data;
  wire [63:0] dcArb_io_requestor_0_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire  dcArb_io_requestor_0_replay_next;
  wire  dcArb_io_requestor_0_xcpt_ma_ld;
  wire  dcArb_io_requestor_0_xcpt_ma_st;
  wire  dcArb_io_requestor_0_xcpt_pf_ld;
  wire  dcArb_io_requestor_0_xcpt_pf_st;
  wire  dcArb_io_requestor_0_invalidate_lr;
  wire  dcArb_io_requestor_0_ordered;
  wire  dcArb_io_mem_req_ready;
  wire  dcArb_io_mem_req_valid;
  wire [39:0] dcArb_io_mem_req_bits_addr;
  wire [5:0] dcArb_io_mem_req_bits_tag;
  wire [4:0] dcArb_io_mem_req_bits_cmd;
  wire [2:0] dcArb_io_mem_req_bits_typ;
  wire  dcArb_io_mem_req_bits_phys;
  wire [63:0] dcArb_io_mem_req_bits_data;
  wire  dcArb_io_mem_s1_kill;
  wire [63:0] dcArb_io_mem_s1_data;
  wire  dcArb_io_mem_s2_nack;
  wire  dcArb_io_mem_resp_valid;
  wire [39:0] dcArb_io_mem_resp_bits_addr;
  wire [5:0] dcArb_io_mem_resp_bits_tag;
  wire [4:0] dcArb_io_mem_resp_bits_cmd;
  wire [2:0] dcArb_io_mem_resp_bits_typ;
  wire [63:0] dcArb_io_mem_resp_bits_data;
  wire  dcArb_io_mem_resp_bits_replay;
  wire  dcArb_io_mem_resp_bits_has_data;
  wire [63:0] dcArb_io_mem_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_mem_resp_bits_store_data;
  wire  dcArb_io_mem_replay_next;
  wire  dcArb_io_mem_xcpt_ma_ld;
  wire  dcArb_io_mem_xcpt_ma_st;
  wire  dcArb_io_mem_xcpt_pf_ld;
  wire  dcArb_io_mem_xcpt_pf_st;
  wire  dcArb_io_mem_invalidate_lr;
  wire  dcArb_io_mem_ordered;
  wire  GEN_0;
  reg [31:0] GEN_160;
  wire [4:0] GEN_1;
  reg [31:0] GEN_161;
  wire [63:0] GEN_2;
  reg [63:0] GEN_162;
  wire [63:0] GEN_3;
  reg [63:0] GEN_163;
  wire  GEN_4;
  reg [31:0] GEN_164;
  wire  GEN_5;
  reg [31:0] GEN_165;
  wire  GEN_6;
  reg [31:0] GEN_166;
  wire [4:0] GEN_7;
  reg [31:0] GEN_167;
  wire  GEN_8;
  reg [31:0] GEN_168;
  wire  GEN_9;
  reg [31:0] GEN_169;
  wire  GEN_10;
  reg [31:0] GEN_170;
  wire  GEN_11;
  reg [31:0] GEN_171;
  wire  GEN_12;
  reg [31:0] GEN_172;
  wire  GEN_13;
  reg [31:0] GEN_173;
  wire  GEN_14;
  reg [31:0] GEN_174;
  wire  GEN_15;
  reg [31:0] GEN_175;
  wire  GEN_16;
  reg [31:0] GEN_176;
  wire  GEN_17;
  reg [31:0] GEN_177;
  wire  GEN_18;
  reg [31:0] GEN_178;
  wire  GEN_19;
  reg [31:0] GEN_179;
  wire  GEN_20;
  reg [31:0] GEN_180;
  wire  GEN_21;
  reg [31:0] GEN_181;
  wire  GEN_22;
  reg [31:0] GEN_182;
  wire  GEN_23;
  reg [31:0] GEN_183;
  wire  GEN_24;
  reg [31:0] GEN_184;
  wire  GEN_25;
  reg [31:0] GEN_185;
  wire [4:0] GEN_26;
  reg [31:0] GEN_186;
  wire  GEN_27;
  reg [31:0] GEN_187;
  wire  GEN_28;
  reg [31:0] GEN_188;
  wire [64:0] GEN_29;
  reg [95:0] GEN_189;
  wire [4:0] GEN_30;
  reg [31:0] GEN_190;
  wire  GEN_31;
  reg [31:0] GEN_191;
  wire  GEN_32;
  reg [31:0] GEN_192;
  wire [4:0] GEN_33;
  reg [31:0] GEN_193;
  wire [63:0] GEN_34;
  reg [63:0] GEN_194;
  wire  GEN_35;
  reg [31:0] GEN_195;
  wire [39:0] GEN_36;
  reg [63:0] GEN_196;
  wire [5:0] GEN_37;
  reg [31:0] GEN_197;
  wire [4:0] GEN_38;
  reg [31:0] GEN_198;
  wire [2:0] GEN_39;
  reg [31:0] GEN_199;
  wire  GEN_40;
  reg [31:0] GEN_200;
  wire [63:0] GEN_41;
  reg [63:0] GEN_201;
  wire  GEN_42;
  reg [31:0] GEN_202;
  wire [63:0] GEN_43;
  reg [63:0] GEN_203;
  wire  GEN_44;
  reg [31:0] GEN_204;
  wire  GEN_45;
  reg [31:0] GEN_205;
  wire  GEN_46;
  reg [31:0] GEN_206;
  wire  GEN_47;
  reg [31:0] GEN_207;
  wire [25:0] GEN_48;
  reg [31:0] GEN_208;
  wire  GEN_49;
  reg [31:0] GEN_209;
  wire [2:0] GEN_50;
  reg [31:0] GEN_210;
  wire  GEN_51;
  reg [31:0] GEN_211;
  wire [2:0] GEN_52;
  reg [31:0] GEN_212;
  wire [10:0] GEN_53;
  reg [31:0] GEN_213;
  wire [63:0] GEN_54;
  reg [63:0] GEN_214;
  wire  GEN_55;
  reg [31:0] GEN_215;
  wire  GEN_56;
  reg [31:0] GEN_216;
  wire [4:0] GEN_57;
  reg [31:0] GEN_217;
  wire  GEN_58;
  reg [31:0] GEN_218;
  wire  GEN_59;
  reg [31:0] GEN_219;
  wire  GEN_60;
  reg [31:0] GEN_220;
  wire  GEN_61;
  reg [31:0] GEN_221;
  wire  GEN_62;
  reg [31:0] GEN_222;
  wire  GEN_63;
  reg [31:0] GEN_223;
  wire  GEN_64;
  reg [31:0] GEN_224;
  wire  GEN_65;
  reg [31:0] GEN_225;
  wire  GEN_66;
  reg [31:0] GEN_226;
  wire  GEN_67;
  reg [31:0] GEN_227;
  wire  GEN_68;
  reg [31:0] GEN_228;
  wire  GEN_69;
  reg [31:0] GEN_229;
  wire  GEN_70;
  reg [31:0] GEN_230;
  wire  GEN_71;
  reg [31:0] GEN_231;
  wire  GEN_72;
  reg [31:0] GEN_232;
  wire  GEN_73;
  reg [31:0] GEN_233;
  wire [2:0] GEN_74;
  reg [31:0] GEN_234;
  wire [1:0] GEN_75;
  reg [31:0] GEN_235;
  wire [64:0] GEN_76;
  reg [95:0] GEN_236;
  wire [64:0] GEN_77;
  reg [95:0] GEN_237;
  wire [64:0] GEN_78;
  reg [95:0] GEN_238;
  wire  GEN_79;
  reg [31:0] GEN_239;
  wire  GEN_80;
  reg [31:0] GEN_240;
  wire  GEN_81;
  reg [31:0] GEN_241;
  wire [15:0] GEN_82;
  reg [31:0] GEN_242;
  wire [37:0] GEN_83;
  reg [63:0] GEN_243;
  wire [1:0] GEN_84;
  reg [31:0] GEN_244;
  wire  GEN_85;
  reg [31:0] GEN_245;
  wire  GEN_86;
  reg [31:0] GEN_246;
  wire  GEN_87;
  reg [31:0] GEN_247;
  wire  GEN_88;
  reg [31:0] GEN_248;
  wire  GEN_89;
  reg [31:0] GEN_249;
  wire  GEN_90;
  reg [31:0] GEN_250;
  wire  GEN_91;
  reg [31:0] GEN_251;
  wire  GEN_92;
  reg [31:0] GEN_252;
  wire [6:0] GEN_93;
  reg [31:0] GEN_253;
  wire [37:0] GEN_94;
  reg [63:0] GEN_254;
  wire  GEN_95;
  reg [31:0] GEN_255;
  wire  GEN_96;
  reg [31:0] GEN_256;
  wire [1:0] GEN_97;
  reg [31:0] GEN_257;
  wire  GEN_98;
  reg [31:0] GEN_258;
  wire [30:0] GEN_99;
  reg [31:0] GEN_259;
  wire  GEN_100;
  reg [31:0] GEN_260;
  wire [1:0] GEN_101;
  reg [31:0] GEN_261;
  wire [4:0] GEN_102;
  reg [31:0] GEN_262;
  wire [3:0] GEN_103;
  reg [31:0] GEN_263;
  wire  GEN_104;
  reg [31:0] GEN_264;
  wire  GEN_105;
  reg [31:0] GEN_265;
  wire  GEN_106;
  reg [31:0] GEN_266;
  wire [1:0] GEN_107;
  reg [31:0] GEN_267;
  wire [1:0] GEN_108;
  reg [31:0] GEN_268;
  wire [1:0] GEN_109;
  reg [31:0] GEN_269;
  wire [1:0] GEN_110;
  reg [31:0] GEN_270;
  wire  GEN_111;
  reg [31:0] GEN_271;
  wire  GEN_112;
  reg [31:0] GEN_272;
  wire  GEN_113;
  reg [31:0] GEN_273;
  wire  GEN_114;
  reg [31:0] GEN_274;
  wire  GEN_115;
  reg [31:0] GEN_275;
  wire  GEN_116;
  reg [31:0] GEN_276;
  wire  GEN_117;
  reg [31:0] GEN_277;
  wire  GEN_118;
  reg [31:0] GEN_278;
  wire  GEN_119;
  reg [31:0] GEN_279;
  wire  GEN_120;
  reg [31:0] GEN_280;
  wire  GEN_121;
  reg [31:0] GEN_281;
  wire [15:0] GEN_122;
  reg [31:0] GEN_282;
  wire [37:0] GEN_123;
  reg [63:0] GEN_283;
  wire [1:0] GEN_124;
  reg [31:0] GEN_284;
  wire  GEN_125;
  reg [31:0] GEN_285;
  wire  GEN_126;
  reg [31:0] GEN_286;
  wire  GEN_127;
  reg [31:0] GEN_287;
  wire  GEN_128;
  reg [31:0] GEN_288;
  wire  GEN_129;
  reg [31:0] GEN_289;
  wire  GEN_130;
  reg [31:0] GEN_290;
  wire  GEN_131;
  reg [31:0] GEN_291;
  wire  GEN_132;
  reg [31:0] GEN_292;
  wire [6:0] GEN_133;
  reg [31:0] GEN_293;
  wire [37:0] GEN_134;
  reg [63:0] GEN_294;
  wire  GEN_135;
  reg [31:0] GEN_295;
  wire  GEN_136;
  reg [31:0] GEN_296;
  wire [1:0] GEN_137;
  reg [31:0] GEN_297;
  wire  GEN_138;
  reg [31:0] GEN_298;
  wire [30:0] GEN_139;
  reg [31:0] GEN_299;
  wire  GEN_140;
  reg [31:0] GEN_300;
  wire [1:0] GEN_141;
  reg [31:0] GEN_301;
  wire [4:0] GEN_142;
  reg [31:0] GEN_302;
  wire [3:0] GEN_143;
  reg [31:0] GEN_303;
  wire  GEN_144;
  reg [31:0] GEN_304;
  wire  GEN_145;
  reg [31:0] GEN_305;
  wire  GEN_146;
  reg [31:0] GEN_306;
  wire [1:0] GEN_147;
  reg [31:0] GEN_307;
  wire [1:0] GEN_148;
  reg [31:0] GEN_308;
  wire [1:0] GEN_149;
  reg [31:0] GEN_309;
  wire [1:0] GEN_150;
  reg [31:0] GEN_310;
  wire  GEN_151;
  reg [31:0] GEN_311;
  wire  GEN_152;
  reg [31:0] GEN_312;
  wire  GEN_153;
  reg [31:0] GEN_313;
  wire  GEN_154;
  reg [31:0] GEN_314;
  wire  GEN_155;
  reg [31:0] GEN_315;
  wire  GEN_156;
  reg [31:0] GEN_316;
  wire  GEN_157;
  reg [31:0] GEN_317;
  wire  GEN_158;
  reg [31:0] GEN_318;
  wire  GEN_159;
  reg [31:0] GEN_319;
  Rocket core (
    .clk(core_clk),
    .reset(core_reset),
    .io_prci_reset(core_io_prci_reset),
    .io_prci_id(core_io_prci_id),
    .io_prci_interrupts_meip(core_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(core_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(core_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(core_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(core_io_prci_interrupts_msip),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_btb_valid(core_io_imem_resp_bits_btb_valid),
    .io_imem_resp_bits_btb_bits_taken(core_io_imem_resp_bits_btb_bits_taken),
    .io_imem_resp_bits_btb_bits_mask(core_io_imem_resp_bits_btb_bits_mask),
    .io_imem_resp_bits_btb_bits_bridx(core_io_imem_resp_bits_btb_bits_bridx),
    .io_imem_resp_bits_btb_bits_target(core_io_imem_resp_bits_btb_bits_target),
    .io_imem_resp_bits_btb_bits_entry(core_io_imem_resp_bits_btb_bits_entry),
    .io_imem_resp_bits_btb_bits_bht_history(core_io_imem_resp_bits_btb_bits_bht_history),
    .io_imem_resp_bits_btb_bits_bht_value(core_io_imem_resp_bits_btb_bits_bht_value),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_imem_resp_bits_mask(core_io_imem_resp_bits_mask),
    .io_imem_resp_bits_xcpt_if(core_io_imem_resp_bits_xcpt_if),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_btb_update_bits_prediction_valid(core_io_imem_btb_update_bits_prediction_valid),
    .io_imem_btb_update_bits_prediction_bits_taken(core_io_imem_btb_update_bits_prediction_bits_taken),
    .io_imem_btb_update_bits_prediction_bits_mask(core_io_imem_btb_update_bits_prediction_bits_mask),
    .io_imem_btb_update_bits_prediction_bits_bridx(core_io_imem_btb_update_bits_prediction_bits_bridx),
    .io_imem_btb_update_bits_prediction_bits_target(core_io_imem_btb_update_bits_prediction_bits_target),
    .io_imem_btb_update_bits_prediction_bits_entry(core_io_imem_btb_update_bits_prediction_bits_entry),
    .io_imem_btb_update_bits_prediction_bits_bht_history(core_io_imem_btb_update_bits_prediction_bits_bht_history),
    .io_imem_btb_update_bits_prediction_bits_bht_value(core_io_imem_btb_update_bits_prediction_bits_bht_value),
    .io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),
    .io_imem_btb_update_bits_target(core_io_imem_btb_update_bits_target),
    .io_imem_btb_update_bits_taken(core_io_imem_btb_update_bits_taken),
    .io_imem_btb_update_bits_isValid(core_io_imem_btb_update_bits_isValid),
    .io_imem_btb_update_bits_isJump(core_io_imem_btb_update_bits_isJump),
    .io_imem_btb_update_bits_isReturn(core_io_imem_btb_update_bits_isReturn),
    .io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_bht_update_bits_prediction_valid(core_io_imem_bht_update_bits_prediction_valid),
    .io_imem_bht_update_bits_prediction_bits_taken(core_io_imem_bht_update_bits_prediction_bits_taken),
    .io_imem_bht_update_bits_prediction_bits_mask(core_io_imem_bht_update_bits_prediction_bits_mask),
    .io_imem_bht_update_bits_prediction_bits_bridx(core_io_imem_bht_update_bits_prediction_bits_bridx),
    .io_imem_bht_update_bits_prediction_bits_target(core_io_imem_bht_update_bits_prediction_bits_target),
    .io_imem_bht_update_bits_prediction_bits_entry(core_io_imem_bht_update_bits_prediction_bits_entry),
    .io_imem_bht_update_bits_prediction_bits_bht_history(core_io_imem_bht_update_bits_prediction_bits_bht_history),
    .io_imem_bht_update_bits_prediction_bits_bht_value(core_io_imem_bht_update_bits_prediction_bits_bht_value),
    .io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),
    .io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),
    .io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),
    .io_imem_ras_update_valid(core_io_imem_ras_update_valid),
    .io_imem_ras_update_bits_isCall(core_io_imem_ras_update_bits_isCall),
    .io_imem_ras_update_bits_isReturn(core_io_imem_ras_update_bits_isReturn),
    .io_imem_ras_update_bits_returnAddr(core_io_imem_ras_update_bits_returnAddr),
    .io_imem_ras_update_bits_prediction_valid(core_io_imem_ras_update_bits_prediction_valid),
    .io_imem_ras_update_bits_prediction_bits_taken(core_io_imem_ras_update_bits_prediction_bits_taken),
    .io_imem_ras_update_bits_prediction_bits_mask(core_io_imem_ras_update_bits_prediction_bits_mask),
    .io_imem_ras_update_bits_prediction_bits_bridx(core_io_imem_ras_update_bits_prediction_bits_bridx),
    .io_imem_ras_update_bits_prediction_bits_target(core_io_imem_ras_update_bits_prediction_bits_target),
    .io_imem_ras_update_bits_prediction_bits_entry(core_io_imem_ras_update_bits_prediction_bits_entry),
    .io_imem_ras_update_bits_prediction_bits_bht_history(core_io_imem_ras_update_bits_prediction_bits_bht_history),
    .io_imem_ras_update_bits_prediction_bits_bht_value(core_io_imem_ras_update_bits_prediction_bits_bht_value),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_imem_flush_tlb(core_io_imem_flush_tlb),
    .io_imem_npc(core_io_imem_npc),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_req_bits_phys(core_io_dmem_req_bits_phys),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data(core_io_dmem_s1_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_addr(core_io_dmem_resp_bits_addr),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_cmd(core_io_dmem_resp_bits_cmd),
    .io_dmem_resp_bits_typ(core_io_dmem_resp_bits_typ),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_resp_bits_store_data(core_io_dmem_resp_bits_store_data),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_xcpt_ma_ld(core_io_dmem_xcpt_ma_ld),
    .io_dmem_xcpt_ma_st(core_io_dmem_xcpt_ma_st),
    .io_dmem_xcpt_pf_ld(core_io_dmem_xcpt_pf_ld),
    .io_dmem_xcpt_pf_st(core_io_dmem_xcpt_pf_st),
    .io_dmem_invalidate_lr(core_io_dmem_invalidate_lr),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_ptw_ptbr_asid(core_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(core_io_ptw_invalidate),
    .io_ptw_status_debug(core_io_ptw_status_debug),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_sd(core_io_ptw_status_sd),
    .io_ptw_status_zero3(core_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(core_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(core_io_ptw_status_zero2),
    .io_ptw_status_vm(core_io_ptw_status_vm),
    .io_ptw_status_zero1(core_io_ptw_status_zero1),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_pum(core_io_ptw_status_pum),
    .io_ptw_status_mprv(core_io_ptw_status_mprv),
    .io_ptw_status_xs(core_io_ptw_status_xs),
    .io_ptw_status_fs(core_io_ptw_status_fs),
    .io_ptw_status_mpp(core_io_ptw_status_mpp),
    .io_ptw_status_hpp(core_io_ptw_status_hpp),
    .io_ptw_status_spp(core_io_ptw_status_spp),
    .io_ptw_status_mpie(core_io_ptw_status_mpie),
    .io_ptw_status_hpie(core_io_ptw_status_hpie),
    .io_ptw_status_spie(core_io_ptw_status_spie),
    .io_ptw_status_upie(core_io_ptw_status_upie),
    .io_ptw_status_mie(core_io_ptw_status_mie),
    .io_ptw_status_hie(core_io_ptw_status_hie),
    .io_ptw_status_sie(core_io_ptw_status_sie),
    .io_ptw_status_uie(core_io_ptw_status_uie),
    .io_fpu_inst(core_io_fpu_inst),
    .io_fpu_fromint_data(core_io_fpu_fromint_data),
    .io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),
    .io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),
    .io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),
    .io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),
    .io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),
    .io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),
    .io_fpu_valid(core_io_fpu_valid),
    .io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_illegal_rm(core_io_fpu_illegal_rm),
    .io_fpu_killx(core_io_fpu_killx),
    .io_fpu_killm(core_io_fpu_killm),
    .io_fpu_dec_cmd(core_io_fpu_dec_cmd),
    .io_fpu_dec_ldst(core_io_fpu_dec_ldst),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_fpu_dec_swap12(core_io_fpu_dec_swap12),
    .io_fpu_dec_swap23(core_io_fpu_dec_swap23),
    .io_fpu_dec_single(core_io_fpu_dec_single),
    .io_fpu_dec_fromint(core_io_fpu_dec_fromint),
    .io_fpu_dec_toint(core_io_fpu_dec_toint),
    .io_fpu_dec_fastpipe(core_io_fpu_dec_fastpipe),
    .io_fpu_dec_fma(core_io_fpu_dec_fma),
    .io_fpu_dec_div(core_io_fpu_dec_div),
    .io_fpu_dec_sqrt(core_io_fpu_dec_sqrt),
    .io_fpu_dec_round(core_io_fpu_dec_round),
    .io_fpu_dec_wflags(core_io_fpu_dec_wflags),
    .io_fpu_sboard_set(core_io_fpu_sboard_set),
    .io_fpu_sboard_clr(core_io_fpu_sboard_clr),
    .io_fpu_sboard_clra(core_io_fpu_sboard_clra),
    .io_fpu_cp_req_ready(core_io_fpu_cp_req_ready),
    .io_fpu_cp_req_valid(core_io_fpu_cp_req_valid),
    .io_fpu_cp_req_bits_cmd(core_io_fpu_cp_req_bits_cmd),
    .io_fpu_cp_req_bits_ldst(core_io_fpu_cp_req_bits_ldst),
    .io_fpu_cp_req_bits_wen(core_io_fpu_cp_req_bits_wen),
    .io_fpu_cp_req_bits_ren1(core_io_fpu_cp_req_bits_ren1),
    .io_fpu_cp_req_bits_ren2(core_io_fpu_cp_req_bits_ren2),
    .io_fpu_cp_req_bits_ren3(core_io_fpu_cp_req_bits_ren3),
    .io_fpu_cp_req_bits_swap12(core_io_fpu_cp_req_bits_swap12),
    .io_fpu_cp_req_bits_swap23(core_io_fpu_cp_req_bits_swap23),
    .io_fpu_cp_req_bits_single(core_io_fpu_cp_req_bits_single),
    .io_fpu_cp_req_bits_fromint(core_io_fpu_cp_req_bits_fromint),
    .io_fpu_cp_req_bits_toint(core_io_fpu_cp_req_bits_toint),
    .io_fpu_cp_req_bits_fastpipe(core_io_fpu_cp_req_bits_fastpipe),
    .io_fpu_cp_req_bits_fma(core_io_fpu_cp_req_bits_fma),
    .io_fpu_cp_req_bits_div(core_io_fpu_cp_req_bits_div),
    .io_fpu_cp_req_bits_sqrt(core_io_fpu_cp_req_bits_sqrt),
    .io_fpu_cp_req_bits_round(core_io_fpu_cp_req_bits_round),
    .io_fpu_cp_req_bits_wflags(core_io_fpu_cp_req_bits_wflags),
    .io_fpu_cp_req_bits_rm(core_io_fpu_cp_req_bits_rm),
    .io_fpu_cp_req_bits_typ(core_io_fpu_cp_req_bits_typ),
    .io_fpu_cp_req_bits_in1(core_io_fpu_cp_req_bits_in1),
    .io_fpu_cp_req_bits_in2(core_io_fpu_cp_req_bits_in2),
    .io_fpu_cp_req_bits_in3(core_io_fpu_cp_req_bits_in3),
    .io_fpu_cp_resp_ready(core_io_fpu_cp_resp_ready),
    .io_fpu_cp_resp_valid(core_io_fpu_cp_resp_valid),
    .io_fpu_cp_resp_bits_data(core_io_fpu_cp_resp_bits_data),
    .io_fpu_cp_resp_bits_exc(core_io_fpu_cp_resp_bits_exc),
    .io_rocc_cmd_ready(core_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(core_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(core_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(core_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(core_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(core_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(core_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(core_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(core_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(core_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(core_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(core_io_rocc_cmd_bits_rs2),
    .io_rocc_cmd_bits_status_debug(core_io_rocc_cmd_bits_status_debug),
    .io_rocc_cmd_bits_status_prv(core_io_rocc_cmd_bits_status_prv),
    .io_rocc_cmd_bits_status_sd(core_io_rocc_cmd_bits_status_sd),
    .io_rocc_cmd_bits_status_zero3(core_io_rocc_cmd_bits_status_zero3),
    .io_rocc_cmd_bits_status_sd_rv32(core_io_rocc_cmd_bits_status_sd_rv32),
    .io_rocc_cmd_bits_status_zero2(core_io_rocc_cmd_bits_status_zero2),
    .io_rocc_cmd_bits_status_vm(core_io_rocc_cmd_bits_status_vm),
    .io_rocc_cmd_bits_status_zero1(core_io_rocc_cmd_bits_status_zero1),
    .io_rocc_cmd_bits_status_mxr(core_io_rocc_cmd_bits_status_mxr),
    .io_rocc_cmd_bits_status_pum(core_io_rocc_cmd_bits_status_pum),
    .io_rocc_cmd_bits_status_mprv(core_io_rocc_cmd_bits_status_mprv),
    .io_rocc_cmd_bits_status_xs(core_io_rocc_cmd_bits_status_xs),
    .io_rocc_cmd_bits_status_fs(core_io_rocc_cmd_bits_status_fs),
    .io_rocc_cmd_bits_status_mpp(core_io_rocc_cmd_bits_status_mpp),
    .io_rocc_cmd_bits_status_hpp(core_io_rocc_cmd_bits_status_hpp),
    .io_rocc_cmd_bits_status_spp(core_io_rocc_cmd_bits_status_spp),
    .io_rocc_cmd_bits_status_mpie(core_io_rocc_cmd_bits_status_mpie),
    .io_rocc_cmd_bits_status_hpie(core_io_rocc_cmd_bits_status_hpie),
    .io_rocc_cmd_bits_status_spie(core_io_rocc_cmd_bits_status_spie),
    .io_rocc_cmd_bits_status_upie(core_io_rocc_cmd_bits_status_upie),
    .io_rocc_cmd_bits_status_mie(core_io_rocc_cmd_bits_status_mie),
    .io_rocc_cmd_bits_status_hie(core_io_rocc_cmd_bits_status_hie),
    .io_rocc_cmd_bits_status_sie(core_io_rocc_cmd_bits_status_sie),
    .io_rocc_cmd_bits_status_uie(core_io_rocc_cmd_bits_status_uie),
    .io_rocc_resp_ready(core_io_rocc_resp_ready),
    .io_rocc_resp_valid(core_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(core_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(core_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(core_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(core_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(core_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(core_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(core_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(core_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(core_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(core_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(core_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(core_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(core_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(core_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(core_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(core_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(core_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(core_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(core_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(core_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(core_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(core_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(core_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(core_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(core_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(core_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(core_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(core_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(core_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(core_io_rocc_mem_ordered),
    .io_rocc_busy(core_io_rocc_busy),
    .io_rocc_interrupt(core_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(core_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(core_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(core_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(core_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(core_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(core_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(core_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(core_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(core_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(core_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(core_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(core_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(core_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(core_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(core_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(core_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(core_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(core_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(core_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(core_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(core_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(core_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(core_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(core_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(core_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(core_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(core_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(core_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(core_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(core_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(core_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(core_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(core_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(core_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(core_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(core_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(core_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(core_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(core_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(core_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(core_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(core_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(core_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(core_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(core_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(core_io_rocc_exception)
  );
  Frontend icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_cpu_req_valid(icache_io_cpu_req_valid),
    .io_cpu_req_bits_pc(icache_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(icache_io_cpu_req_bits_speculative),
    .io_cpu_resp_ready(icache_io_cpu_resp_ready),
    .io_cpu_resp_valid(icache_io_cpu_resp_valid),
    .io_cpu_resp_bits_btb_valid(icache_io_cpu_resp_bits_btb_valid),
    .io_cpu_resp_bits_btb_bits_taken(icache_io_cpu_resp_bits_btb_bits_taken),
    .io_cpu_resp_bits_btb_bits_mask(icache_io_cpu_resp_bits_btb_bits_mask),
    .io_cpu_resp_bits_btb_bits_bridx(icache_io_cpu_resp_bits_btb_bits_bridx),
    .io_cpu_resp_bits_btb_bits_target(icache_io_cpu_resp_bits_btb_bits_target),
    .io_cpu_resp_bits_btb_bits_entry(icache_io_cpu_resp_bits_btb_bits_entry),
    .io_cpu_resp_bits_btb_bits_bht_history(icache_io_cpu_resp_bits_btb_bits_bht_history),
    .io_cpu_resp_bits_btb_bits_bht_value(icache_io_cpu_resp_bits_btb_bits_bht_value),
    .io_cpu_resp_bits_pc(icache_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data(icache_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_mask(icache_io_cpu_resp_bits_mask),
    .io_cpu_resp_bits_xcpt_if(icache_io_cpu_resp_bits_xcpt_if),
    .io_cpu_resp_bits_replay(icache_io_cpu_resp_bits_replay),
    .io_cpu_btb_update_valid(icache_io_cpu_btb_update_valid),
    .io_cpu_btb_update_bits_prediction_valid(icache_io_cpu_btb_update_bits_prediction_valid),
    .io_cpu_btb_update_bits_prediction_bits_taken(icache_io_cpu_btb_update_bits_prediction_bits_taken),
    .io_cpu_btb_update_bits_prediction_bits_mask(icache_io_cpu_btb_update_bits_prediction_bits_mask),
    .io_cpu_btb_update_bits_prediction_bits_bridx(icache_io_cpu_btb_update_bits_prediction_bits_bridx),
    .io_cpu_btb_update_bits_prediction_bits_target(icache_io_cpu_btb_update_bits_prediction_bits_target),
    .io_cpu_btb_update_bits_prediction_bits_entry(icache_io_cpu_btb_update_bits_prediction_bits_entry),
    .io_cpu_btb_update_bits_prediction_bits_bht_history(icache_io_cpu_btb_update_bits_prediction_bits_bht_history),
    .io_cpu_btb_update_bits_prediction_bits_bht_value(icache_io_cpu_btb_update_bits_prediction_bits_bht_value),
    .io_cpu_btb_update_bits_pc(icache_io_cpu_btb_update_bits_pc),
    .io_cpu_btb_update_bits_target(icache_io_cpu_btb_update_bits_target),
    .io_cpu_btb_update_bits_taken(icache_io_cpu_btb_update_bits_taken),
    .io_cpu_btb_update_bits_isValid(icache_io_cpu_btb_update_bits_isValid),
    .io_cpu_btb_update_bits_isJump(icache_io_cpu_btb_update_bits_isJump),
    .io_cpu_btb_update_bits_isReturn(icache_io_cpu_btb_update_bits_isReturn),
    .io_cpu_btb_update_bits_br_pc(icache_io_cpu_btb_update_bits_br_pc),
    .io_cpu_bht_update_valid(icache_io_cpu_bht_update_valid),
    .io_cpu_bht_update_bits_prediction_valid(icache_io_cpu_bht_update_bits_prediction_valid),
    .io_cpu_bht_update_bits_prediction_bits_taken(icache_io_cpu_bht_update_bits_prediction_bits_taken),
    .io_cpu_bht_update_bits_prediction_bits_mask(icache_io_cpu_bht_update_bits_prediction_bits_mask),
    .io_cpu_bht_update_bits_prediction_bits_bridx(icache_io_cpu_bht_update_bits_prediction_bits_bridx),
    .io_cpu_bht_update_bits_prediction_bits_target(icache_io_cpu_bht_update_bits_prediction_bits_target),
    .io_cpu_bht_update_bits_prediction_bits_entry(icache_io_cpu_bht_update_bits_prediction_bits_entry),
    .io_cpu_bht_update_bits_prediction_bits_bht_history(icache_io_cpu_bht_update_bits_prediction_bits_bht_history),
    .io_cpu_bht_update_bits_prediction_bits_bht_value(icache_io_cpu_bht_update_bits_prediction_bits_bht_value),
    .io_cpu_bht_update_bits_pc(icache_io_cpu_bht_update_bits_pc),
    .io_cpu_bht_update_bits_taken(icache_io_cpu_bht_update_bits_taken),
    .io_cpu_bht_update_bits_mispredict(icache_io_cpu_bht_update_bits_mispredict),
    .io_cpu_ras_update_valid(icache_io_cpu_ras_update_valid),
    .io_cpu_ras_update_bits_isCall(icache_io_cpu_ras_update_bits_isCall),
    .io_cpu_ras_update_bits_isReturn(icache_io_cpu_ras_update_bits_isReturn),
    .io_cpu_ras_update_bits_returnAddr(icache_io_cpu_ras_update_bits_returnAddr),
    .io_cpu_ras_update_bits_prediction_valid(icache_io_cpu_ras_update_bits_prediction_valid),
    .io_cpu_ras_update_bits_prediction_bits_taken(icache_io_cpu_ras_update_bits_prediction_bits_taken),
    .io_cpu_ras_update_bits_prediction_bits_mask(icache_io_cpu_ras_update_bits_prediction_bits_mask),
    .io_cpu_ras_update_bits_prediction_bits_bridx(icache_io_cpu_ras_update_bits_prediction_bits_bridx),
    .io_cpu_ras_update_bits_prediction_bits_target(icache_io_cpu_ras_update_bits_prediction_bits_target),
    .io_cpu_ras_update_bits_prediction_bits_entry(icache_io_cpu_ras_update_bits_prediction_bits_entry),
    .io_cpu_ras_update_bits_prediction_bits_bht_history(icache_io_cpu_ras_update_bits_prediction_bits_bht_history),
    .io_cpu_ras_update_bits_prediction_bits_bht_value(icache_io_cpu_ras_update_bits_prediction_bits_bht_value),
    .io_cpu_flush_icache(icache_io_cpu_flush_icache),
    .io_cpu_flush_tlb(icache_io_cpu_flush_tlb),
    .io_cpu_npc(icache_io_cpu_npc),
    .io_ptw_req_ready(icache_io_ptw_req_ready),
    .io_ptw_req_valid(icache_io_ptw_req_valid),
    .io_ptw_req_bits_prv(icache_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(icache_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(icache_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(icache_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(icache_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(icache_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(icache_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(icache_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(icache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(icache_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(icache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(icache_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(icache_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(icache_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(icache_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(icache_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(icache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(icache_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(icache_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(icache_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(icache_io_ptw_invalidate),
    .io_ptw_status_debug(icache_io_ptw_status_debug),
    .io_ptw_status_prv(icache_io_ptw_status_prv),
    .io_ptw_status_sd(icache_io_ptw_status_sd),
    .io_ptw_status_zero3(icache_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(icache_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(icache_io_ptw_status_zero2),
    .io_ptw_status_vm(icache_io_ptw_status_vm),
    .io_ptw_status_zero1(icache_io_ptw_status_zero1),
    .io_ptw_status_mxr(icache_io_ptw_status_mxr),
    .io_ptw_status_pum(icache_io_ptw_status_pum),
    .io_ptw_status_mprv(icache_io_ptw_status_mprv),
    .io_ptw_status_xs(icache_io_ptw_status_xs),
    .io_ptw_status_fs(icache_io_ptw_status_fs),
    .io_ptw_status_mpp(icache_io_ptw_status_mpp),
    .io_ptw_status_hpp(icache_io_ptw_status_hpp),
    .io_ptw_status_spp(icache_io_ptw_status_spp),
    .io_ptw_status_mpie(icache_io_ptw_status_mpie),
    .io_ptw_status_hpie(icache_io_ptw_status_hpie),
    .io_ptw_status_spie(icache_io_ptw_status_spie),
    .io_ptw_status_upie(icache_io_ptw_status_upie),
    .io_ptw_status_mie(icache_io_ptw_status_mie),
    .io_ptw_status_hie(icache_io_ptw_status_hie),
    .io_ptw_status_sie(icache_io_ptw_status_sie),
    .io_ptw_status_uie(icache_io_ptw_status_uie),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  DCache DCache_1 (
    .clk(DCache_1_clk),
    .reset(DCache_1_reset),
    .io_cpu_req_ready(DCache_1_io_cpu_req_ready),
    .io_cpu_req_valid(DCache_1_io_cpu_req_valid),
    .io_cpu_req_bits_addr(DCache_1_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(DCache_1_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(DCache_1_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_typ(DCache_1_io_cpu_req_bits_typ),
    .io_cpu_req_bits_phys(DCache_1_io_cpu_req_bits_phys),
    .io_cpu_req_bits_data(DCache_1_io_cpu_req_bits_data),
    .io_cpu_s1_kill(DCache_1_io_cpu_s1_kill),
    .io_cpu_s1_data(DCache_1_io_cpu_s1_data),
    .io_cpu_s2_nack(DCache_1_io_cpu_s2_nack),
    .io_cpu_resp_valid(DCache_1_io_cpu_resp_valid),
    .io_cpu_resp_bits_addr(DCache_1_io_cpu_resp_bits_addr),
    .io_cpu_resp_bits_tag(DCache_1_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_cmd(DCache_1_io_cpu_resp_bits_cmd),
    .io_cpu_resp_bits_typ(DCache_1_io_cpu_resp_bits_typ),
    .io_cpu_resp_bits_data(DCache_1_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(DCache_1_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(DCache_1_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(DCache_1_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_resp_bits_store_data(DCache_1_io_cpu_resp_bits_store_data),
    .io_cpu_replay_next(DCache_1_io_cpu_replay_next),
    .io_cpu_xcpt_ma_ld(DCache_1_io_cpu_xcpt_ma_ld),
    .io_cpu_xcpt_ma_st(DCache_1_io_cpu_xcpt_ma_st),
    .io_cpu_xcpt_pf_ld(DCache_1_io_cpu_xcpt_pf_ld),
    .io_cpu_xcpt_pf_st(DCache_1_io_cpu_xcpt_pf_st),
    .io_cpu_invalidate_lr(DCache_1_io_cpu_invalidate_lr),
    .io_cpu_ordered(DCache_1_io_cpu_ordered),
    .io_ptw_req_ready(DCache_1_io_ptw_req_ready),
    .io_ptw_req_valid(DCache_1_io_ptw_req_valid),
    .io_ptw_req_bits_prv(DCache_1_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(DCache_1_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(DCache_1_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(DCache_1_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(DCache_1_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(DCache_1_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(DCache_1_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(DCache_1_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(DCache_1_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(DCache_1_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(DCache_1_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(DCache_1_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(DCache_1_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(DCache_1_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(DCache_1_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(DCache_1_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(DCache_1_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(DCache_1_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(DCache_1_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(DCache_1_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(DCache_1_io_ptw_invalidate),
    .io_ptw_status_debug(DCache_1_io_ptw_status_debug),
    .io_ptw_status_prv(DCache_1_io_ptw_status_prv),
    .io_ptw_status_sd(DCache_1_io_ptw_status_sd),
    .io_ptw_status_zero3(DCache_1_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(DCache_1_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(DCache_1_io_ptw_status_zero2),
    .io_ptw_status_vm(DCache_1_io_ptw_status_vm),
    .io_ptw_status_zero1(DCache_1_io_ptw_status_zero1),
    .io_ptw_status_mxr(DCache_1_io_ptw_status_mxr),
    .io_ptw_status_pum(DCache_1_io_ptw_status_pum),
    .io_ptw_status_mprv(DCache_1_io_ptw_status_mprv),
    .io_ptw_status_xs(DCache_1_io_ptw_status_xs),
    .io_ptw_status_fs(DCache_1_io_ptw_status_fs),
    .io_ptw_status_mpp(DCache_1_io_ptw_status_mpp),
    .io_ptw_status_hpp(DCache_1_io_ptw_status_hpp),
    .io_ptw_status_spp(DCache_1_io_ptw_status_spp),
    .io_ptw_status_mpie(DCache_1_io_ptw_status_mpie),
    .io_ptw_status_hpie(DCache_1_io_ptw_status_hpie),
    .io_ptw_status_spie(DCache_1_io_ptw_status_spie),
    .io_ptw_status_upie(DCache_1_io_ptw_status_upie),
    .io_ptw_status_mie(DCache_1_io_ptw_status_mie),
    .io_ptw_status_hie(DCache_1_io_ptw_status_hie),
    .io_ptw_status_sie(DCache_1_io_ptw_status_sie),
    .io_ptw_status_uie(DCache_1_io_ptw_status_uie),
    .io_mem_acquire_ready(DCache_1_io_mem_acquire_ready),
    .io_mem_acquire_valid(DCache_1_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(DCache_1_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(DCache_1_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(DCache_1_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(DCache_1_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(DCache_1_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(DCache_1_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(DCache_1_io_mem_acquire_bits_data),
    .io_mem_probe_ready(DCache_1_io_mem_probe_ready),
    .io_mem_probe_valid(DCache_1_io_mem_probe_valid),
    .io_mem_probe_bits_addr_block(DCache_1_io_mem_probe_bits_addr_block),
    .io_mem_probe_bits_p_type(DCache_1_io_mem_probe_bits_p_type),
    .io_mem_release_ready(DCache_1_io_mem_release_ready),
    .io_mem_release_valid(DCache_1_io_mem_release_valid),
    .io_mem_release_bits_addr_beat(DCache_1_io_mem_release_bits_addr_beat),
    .io_mem_release_bits_addr_block(DCache_1_io_mem_release_bits_addr_block),
    .io_mem_release_bits_client_xact_id(DCache_1_io_mem_release_bits_client_xact_id),
    .io_mem_release_bits_voluntary(DCache_1_io_mem_release_bits_voluntary),
    .io_mem_release_bits_r_type(DCache_1_io_mem_release_bits_r_type),
    .io_mem_release_bits_data(DCache_1_io_mem_release_bits_data),
    .io_mem_grant_ready(DCache_1_io_mem_grant_ready),
    .io_mem_grant_valid(DCache_1_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(DCache_1_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(DCache_1_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(DCache_1_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(DCache_1_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(DCache_1_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(DCache_1_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(DCache_1_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(DCache_1_io_mem_finish_ready),
    .io_mem_finish_valid(DCache_1_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(DCache_1_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(DCache_1_io_mem_finish_bits_manager_id)
  );
  ClientUncachedTileLinkIOArbiter uncachedArb (
    .clk(uncachedArb_clk),
    .reset(uncachedArb_reset),
    .io_in_0_acquire_ready(uncachedArb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(uncachedArb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(uncachedArb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(uncachedArb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(uncachedArb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(uncachedArb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(uncachedArb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(uncachedArb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(uncachedArb_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(uncachedArb_io_in_0_grant_ready),
    .io_in_0_grant_valid(uncachedArb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(uncachedArb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(uncachedArb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(uncachedArb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(uncachedArb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(uncachedArb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(uncachedArb_io_in_0_grant_bits_data),
    .io_out_acquire_ready(uncachedArb_io_out_acquire_ready),
    .io_out_acquire_valid(uncachedArb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(uncachedArb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(uncachedArb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(uncachedArb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(uncachedArb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(uncachedArb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(uncachedArb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(uncachedArb_io_out_acquire_bits_data),
    .io_out_grant_ready(uncachedArb_io_out_grant_ready),
    .io_out_grant_valid(uncachedArb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(uncachedArb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(uncachedArb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(uncachedArb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(uncachedArb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(uncachedArb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(uncachedArb_io_out_grant_bits_data)
  );
  HellaCacheArbiter dcArb (
    .clk(dcArb_clk),
    .reset(dcArb_reset),
    .io_requestor_0_req_ready(dcArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_tag(dcArb_io_requestor_0_req_bits_tag),
    .io_requestor_0_req_bits_cmd(dcArb_io_requestor_0_req_bits_cmd),
    .io_requestor_0_req_bits_typ(dcArb_io_requestor_0_req_bits_typ),
    .io_requestor_0_req_bits_phys(dcArb_io_requestor_0_req_bits_phys),
    .io_requestor_0_req_bits_data(dcArb_io_requestor_0_req_bits_data),
    .io_requestor_0_s1_kill(dcArb_io_requestor_0_s1_kill),
    .io_requestor_0_s1_data(dcArb_io_requestor_0_s1_data),
    .io_requestor_0_s2_nack(dcArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_addr(dcArb_io_requestor_0_resp_bits_addr),
    .io_requestor_0_resp_bits_tag(dcArb_io_requestor_0_resp_bits_tag),
    .io_requestor_0_resp_bits_cmd(dcArb_io_requestor_0_resp_bits_cmd),
    .io_requestor_0_resp_bits_typ(dcArb_io_requestor_0_resp_bits_typ),
    .io_requestor_0_resp_bits_data(dcArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_resp_bits_replay(dcArb_io_requestor_0_resp_bits_replay),
    .io_requestor_0_resp_bits_has_data(dcArb_io_requestor_0_resp_bits_has_data),
    .io_requestor_0_resp_bits_data_word_bypass(dcArb_io_requestor_0_resp_bits_data_word_bypass),
    .io_requestor_0_resp_bits_store_data(dcArb_io_requestor_0_resp_bits_store_data),
    .io_requestor_0_replay_next(dcArb_io_requestor_0_replay_next),
    .io_requestor_0_xcpt_ma_ld(dcArb_io_requestor_0_xcpt_ma_ld),
    .io_requestor_0_xcpt_ma_st(dcArb_io_requestor_0_xcpt_ma_st),
    .io_requestor_0_xcpt_pf_ld(dcArb_io_requestor_0_xcpt_pf_ld),
    .io_requestor_0_xcpt_pf_st(dcArb_io_requestor_0_xcpt_pf_st),
    .io_requestor_0_invalidate_lr(dcArb_io_requestor_0_invalidate_lr),
    .io_requestor_0_ordered(dcArb_io_requestor_0_ordered),
    .io_mem_req_ready(dcArb_io_mem_req_ready),
    .io_mem_req_valid(dcArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(dcArb_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(dcArb_io_mem_req_bits_phys),
    .io_mem_req_bits_data(dcArb_io_mem_req_bits_data),
    .io_mem_s1_kill(dcArb_io_mem_s1_kill),
    .io_mem_s1_data(dcArb_io_mem_s1_data),
    .io_mem_s2_nack(dcArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcArb_io_mem_resp_valid),
    .io_mem_resp_bits_addr(dcArb_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(dcArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(dcArb_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_typ(dcArb_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(dcArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_store_data(dcArb_io_mem_resp_bits_store_data),
    .io_mem_replay_next(dcArb_io_mem_replay_next),
    .io_mem_xcpt_ma_ld(dcArb_io_mem_xcpt_ma_ld),
    .io_mem_xcpt_ma_st(dcArb_io_mem_xcpt_ma_st),
    .io_mem_xcpt_pf_ld(dcArb_io_mem_xcpt_pf_ld),
    .io_mem_xcpt_pf_st(dcArb_io_mem_xcpt_pf_st),
    .io_mem_invalidate_lr(dcArb_io_mem_invalidate_lr),
    .io_mem_ordered(dcArb_io_mem_ordered)
  );
  assign io_cached_0_acquire_valid = DCache_1_io_mem_acquire_valid;
  assign io_cached_0_acquire_bits_addr_block = DCache_1_io_mem_acquire_bits_addr_block;
  assign io_cached_0_acquire_bits_client_xact_id = DCache_1_io_mem_acquire_bits_client_xact_id;
  assign io_cached_0_acquire_bits_addr_beat = DCache_1_io_mem_acquire_bits_addr_beat;
  assign io_cached_0_acquire_bits_is_builtin_type = DCache_1_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_0_acquire_bits_a_type = DCache_1_io_mem_acquire_bits_a_type;
  assign io_cached_0_acquire_bits_union = DCache_1_io_mem_acquire_bits_union;
  assign io_cached_0_acquire_bits_data = DCache_1_io_mem_acquire_bits_data;
  assign io_cached_0_probe_ready = DCache_1_io_mem_probe_ready;
  assign io_cached_0_release_valid = DCache_1_io_mem_release_valid;
  assign io_cached_0_release_bits_addr_beat = DCache_1_io_mem_release_bits_addr_beat;
  assign io_cached_0_release_bits_addr_block = DCache_1_io_mem_release_bits_addr_block;
  assign io_cached_0_release_bits_client_xact_id = DCache_1_io_mem_release_bits_client_xact_id;
  assign io_cached_0_release_bits_voluntary = DCache_1_io_mem_release_bits_voluntary;
  assign io_cached_0_release_bits_r_type = DCache_1_io_mem_release_bits_r_type;
  assign io_cached_0_release_bits_data = DCache_1_io_mem_release_bits_data;
  assign io_cached_0_grant_ready = DCache_1_io_mem_grant_ready;
  assign io_cached_0_finish_valid = DCache_1_io_mem_finish_valid;
  assign io_cached_0_finish_bits_manager_xact_id = DCache_1_io_mem_finish_bits_manager_xact_id;
  assign io_cached_0_finish_bits_manager_id = DCache_1_io_mem_finish_bits_manager_id;
  assign io_uncached_0_acquire_valid = uncachedArb_io_out_acquire_valid;
  assign io_uncached_0_acquire_bits_addr_block = uncachedArb_io_out_acquire_bits_addr_block;
  assign io_uncached_0_acquire_bits_client_xact_id = uncachedArb_io_out_acquire_bits_client_xact_id;
  assign io_uncached_0_acquire_bits_addr_beat = uncachedArb_io_out_acquire_bits_addr_beat;
  assign io_uncached_0_acquire_bits_is_builtin_type = uncachedArb_io_out_acquire_bits_is_builtin_type;
  assign io_uncached_0_acquire_bits_a_type = uncachedArb_io_out_acquire_bits_a_type;
  assign io_uncached_0_acquire_bits_union = uncachedArb_io_out_acquire_bits_union;
  assign io_uncached_0_acquire_bits_data = uncachedArb_io_out_acquire_bits_data;
  assign io_uncached_0_grant_ready = uncachedArb_io_out_grant_ready;
  assign core_clk = clk;
  assign core_reset = reset;
  assign core_io_prci_reset = io_prci_reset;
  assign core_io_prci_id = io_prci_id;
  assign core_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign core_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign core_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign core_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign core_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign core_io_imem_resp_valid = icache_io_cpu_resp_valid;
  assign core_io_imem_resp_bits_btb_valid = icache_io_cpu_resp_bits_btb_valid;
  assign core_io_imem_resp_bits_btb_bits_taken = icache_io_cpu_resp_bits_btb_bits_taken;
  assign core_io_imem_resp_bits_btb_bits_mask = icache_io_cpu_resp_bits_btb_bits_mask;
  assign core_io_imem_resp_bits_btb_bits_bridx = icache_io_cpu_resp_bits_btb_bits_bridx;
  assign core_io_imem_resp_bits_btb_bits_target = icache_io_cpu_resp_bits_btb_bits_target;
  assign core_io_imem_resp_bits_btb_bits_entry = icache_io_cpu_resp_bits_btb_bits_entry;
  assign core_io_imem_resp_bits_btb_bits_bht_history = icache_io_cpu_resp_bits_btb_bits_bht_history;
  assign core_io_imem_resp_bits_btb_bits_bht_value = icache_io_cpu_resp_bits_btb_bits_bht_value;
  assign core_io_imem_resp_bits_pc = icache_io_cpu_resp_bits_pc;
  assign core_io_imem_resp_bits_data = icache_io_cpu_resp_bits_data;
  assign core_io_imem_resp_bits_mask = icache_io_cpu_resp_bits_mask;
  assign core_io_imem_resp_bits_xcpt_if = icache_io_cpu_resp_bits_xcpt_if;
  assign core_io_imem_resp_bits_replay = icache_io_cpu_resp_bits_replay;
  assign core_io_imem_npc = icache_io_cpu_npc;
  assign core_io_dmem_req_ready = dcArb_io_requestor_0_req_ready;
  assign core_io_dmem_s2_nack = dcArb_io_requestor_0_s2_nack;
  assign core_io_dmem_resp_valid = dcArb_io_requestor_0_resp_valid;
  assign core_io_dmem_resp_bits_addr = dcArb_io_requestor_0_resp_bits_addr;
  assign core_io_dmem_resp_bits_tag = dcArb_io_requestor_0_resp_bits_tag;
  assign core_io_dmem_resp_bits_cmd = dcArb_io_requestor_0_resp_bits_cmd;
  assign core_io_dmem_resp_bits_typ = dcArb_io_requestor_0_resp_bits_typ;
  assign core_io_dmem_resp_bits_data = dcArb_io_requestor_0_resp_bits_data;
  assign core_io_dmem_resp_bits_replay = dcArb_io_requestor_0_resp_bits_replay;
  assign core_io_dmem_resp_bits_has_data = dcArb_io_requestor_0_resp_bits_has_data;
  assign core_io_dmem_resp_bits_data_word_bypass = dcArb_io_requestor_0_resp_bits_data_word_bypass;
  assign core_io_dmem_resp_bits_store_data = dcArb_io_requestor_0_resp_bits_store_data;
  assign core_io_dmem_replay_next = dcArb_io_requestor_0_replay_next;
  assign core_io_dmem_xcpt_ma_ld = dcArb_io_requestor_0_xcpt_ma_ld;
  assign core_io_dmem_xcpt_ma_st = dcArb_io_requestor_0_xcpt_ma_st;
  assign core_io_dmem_xcpt_pf_ld = dcArb_io_requestor_0_xcpt_pf_ld;
  assign core_io_dmem_xcpt_pf_st = dcArb_io_requestor_0_xcpt_pf_st;
  assign core_io_dmem_ordered = dcArb_io_requestor_0_ordered;
  assign core_io_fpu_fcsr_flags_valid = GEN_0;
  assign core_io_fpu_fcsr_flags_bits = GEN_1;
  assign core_io_fpu_store_data = GEN_2;
  assign core_io_fpu_toint_data = GEN_3;
  assign core_io_fpu_fcsr_rdy = GEN_4;
  assign core_io_fpu_nack_mem = GEN_5;
  assign core_io_fpu_illegal_rm = GEN_6;
  assign core_io_fpu_dec_cmd = GEN_7;
  assign core_io_fpu_dec_ldst = GEN_8;
  assign core_io_fpu_dec_wen = GEN_9;
  assign core_io_fpu_dec_ren1 = GEN_10;
  assign core_io_fpu_dec_ren2 = GEN_11;
  assign core_io_fpu_dec_ren3 = GEN_12;
  assign core_io_fpu_dec_swap12 = GEN_13;
  assign core_io_fpu_dec_swap23 = GEN_14;
  assign core_io_fpu_dec_single = GEN_15;
  assign core_io_fpu_dec_fromint = GEN_16;
  assign core_io_fpu_dec_toint = GEN_17;
  assign core_io_fpu_dec_fastpipe = GEN_18;
  assign core_io_fpu_dec_fma = GEN_19;
  assign core_io_fpu_dec_div = GEN_20;
  assign core_io_fpu_dec_sqrt = GEN_21;
  assign core_io_fpu_dec_round = GEN_22;
  assign core_io_fpu_dec_wflags = GEN_23;
  assign core_io_fpu_sboard_set = GEN_24;
  assign core_io_fpu_sboard_clr = GEN_25;
  assign core_io_fpu_sboard_clra = GEN_26;
  assign core_io_fpu_cp_req_ready = GEN_27;
  assign core_io_fpu_cp_resp_valid = GEN_28;
  assign core_io_fpu_cp_resp_bits_data = GEN_29;
  assign core_io_fpu_cp_resp_bits_exc = GEN_30;
  assign core_io_rocc_cmd_ready = GEN_31;
  assign core_io_rocc_resp_valid = GEN_32;
  assign core_io_rocc_resp_bits_rd = GEN_33;
  assign core_io_rocc_resp_bits_data = GEN_34;
  assign core_io_rocc_mem_req_valid = GEN_35;
  assign core_io_rocc_mem_req_bits_addr = GEN_36;
  assign core_io_rocc_mem_req_bits_tag = GEN_37;
  assign core_io_rocc_mem_req_bits_cmd = GEN_38;
  assign core_io_rocc_mem_req_bits_typ = GEN_39;
  assign core_io_rocc_mem_req_bits_phys = GEN_40;
  assign core_io_rocc_mem_req_bits_data = GEN_41;
  assign core_io_rocc_mem_s1_kill = GEN_42;
  assign core_io_rocc_mem_s1_data = GEN_43;
  assign core_io_rocc_mem_invalidate_lr = GEN_44;
  assign core_io_rocc_busy = GEN_45;
  assign core_io_rocc_interrupt = GEN_46;
  assign core_io_rocc_autl_acquire_valid = GEN_47;
  assign core_io_rocc_autl_acquire_bits_addr_block = GEN_48;
  assign core_io_rocc_autl_acquire_bits_client_xact_id = GEN_49;
  assign core_io_rocc_autl_acquire_bits_addr_beat = GEN_50;
  assign core_io_rocc_autl_acquire_bits_is_builtin_type = GEN_51;
  assign core_io_rocc_autl_acquire_bits_a_type = GEN_52;
  assign core_io_rocc_autl_acquire_bits_union = GEN_53;
  assign core_io_rocc_autl_acquire_bits_data = GEN_54;
  assign core_io_rocc_autl_grant_ready = GEN_55;
  assign core_io_rocc_fpu_req_valid = GEN_56;
  assign core_io_rocc_fpu_req_bits_cmd = GEN_57;
  assign core_io_rocc_fpu_req_bits_ldst = GEN_58;
  assign core_io_rocc_fpu_req_bits_wen = GEN_59;
  assign core_io_rocc_fpu_req_bits_ren1 = GEN_60;
  assign core_io_rocc_fpu_req_bits_ren2 = GEN_61;
  assign core_io_rocc_fpu_req_bits_ren3 = GEN_62;
  assign core_io_rocc_fpu_req_bits_swap12 = GEN_63;
  assign core_io_rocc_fpu_req_bits_swap23 = GEN_64;
  assign core_io_rocc_fpu_req_bits_single = GEN_65;
  assign core_io_rocc_fpu_req_bits_fromint = GEN_66;
  assign core_io_rocc_fpu_req_bits_toint = GEN_67;
  assign core_io_rocc_fpu_req_bits_fastpipe = GEN_68;
  assign core_io_rocc_fpu_req_bits_fma = GEN_69;
  assign core_io_rocc_fpu_req_bits_div = GEN_70;
  assign core_io_rocc_fpu_req_bits_sqrt = GEN_71;
  assign core_io_rocc_fpu_req_bits_round = GEN_72;
  assign core_io_rocc_fpu_req_bits_wflags = GEN_73;
  assign core_io_rocc_fpu_req_bits_rm = GEN_74;
  assign core_io_rocc_fpu_req_bits_typ = GEN_75;
  assign core_io_rocc_fpu_req_bits_in1 = GEN_76;
  assign core_io_rocc_fpu_req_bits_in2 = GEN_77;
  assign core_io_rocc_fpu_req_bits_in3 = GEN_78;
  assign core_io_rocc_fpu_resp_ready = GEN_79;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_cpu_req_valid = core_io_imem_req_valid;
  assign icache_io_cpu_req_bits_pc = core_io_imem_req_bits_pc;
  assign icache_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative;
  assign icache_io_cpu_resp_ready = core_io_imem_resp_ready;
  assign icache_io_cpu_btb_update_valid = core_io_imem_btb_update_valid;
  assign icache_io_cpu_btb_update_bits_prediction_valid = core_io_imem_btb_update_bits_prediction_valid;
  assign icache_io_cpu_btb_update_bits_prediction_bits_taken = core_io_imem_btb_update_bits_prediction_bits_taken;
  assign icache_io_cpu_btb_update_bits_prediction_bits_mask = core_io_imem_btb_update_bits_prediction_bits_mask;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bridx = core_io_imem_btb_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_btb_update_bits_prediction_bits_target = core_io_imem_btb_update_bits_prediction_bits_target;
  assign icache_io_cpu_btb_update_bits_prediction_bits_entry = core_io_imem_btb_update_bits_prediction_bits_entry;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_history = core_io_imem_btb_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_value = core_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_btb_update_bits_pc = core_io_imem_btb_update_bits_pc;
  assign icache_io_cpu_btb_update_bits_target = core_io_imem_btb_update_bits_target;
  assign icache_io_cpu_btb_update_bits_taken = core_io_imem_btb_update_bits_taken;
  assign icache_io_cpu_btb_update_bits_isValid = core_io_imem_btb_update_bits_isValid;
  assign icache_io_cpu_btb_update_bits_isJump = core_io_imem_btb_update_bits_isJump;
  assign icache_io_cpu_btb_update_bits_isReturn = core_io_imem_btb_update_bits_isReturn;
  assign icache_io_cpu_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc;
  assign icache_io_cpu_bht_update_valid = core_io_imem_bht_update_valid;
  assign icache_io_cpu_bht_update_bits_prediction_valid = core_io_imem_bht_update_bits_prediction_valid;
  assign icache_io_cpu_bht_update_bits_prediction_bits_taken = core_io_imem_bht_update_bits_prediction_bits_taken;
  assign icache_io_cpu_bht_update_bits_prediction_bits_mask = core_io_imem_bht_update_bits_prediction_bits_mask;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bridx = core_io_imem_bht_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_bht_update_bits_prediction_bits_target = core_io_imem_bht_update_bits_prediction_bits_target;
  assign icache_io_cpu_bht_update_bits_prediction_bits_entry = core_io_imem_bht_update_bits_prediction_bits_entry;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_history = core_io_imem_bht_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_value = core_io_imem_bht_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_bht_update_bits_pc = core_io_imem_bht_update_bits_pc;
  assign icache_io_cpu_bht_update_bits_taken = core_io_imem_bht_update_bits_taken;
  assign icache_io_cpu_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict;
  assign icache_io_cpu_ras_update_valid = core_io_imem_ras_update_valid;
  assign icache_io_cpu_ras_update_bits_isCall = core_io_imem_ras_update_bits_isCall;
  assign icache_io_cpu_ras_update_bits_isReturn = core_io_imem_ras_update_bits_isReturn;
  assign icache_io_cpu_ras_update_bits_returnAddr = core_io_imem_ras_update_bits_returnAddr;
  assign icache_io_cpu_ras_update_bits_prediction_valid = core_io_imem_ras_update_bits_prediction_valid;
  assign icache_io_cpu_ras_update_bits_prediction_bits_taken = core_io_imem_ras_update_bits_prediction_bits_taken;
  assign icache_io_cpu_ras_update_bits_prediction_bits_mask = core_io_imem_ras_update_bits_prediction_bits_mask;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bridx = core_io_imem_ras_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_ras_update_bits_prediction_bits_target = core_io_imem_ras_update_bits_prediction_bits_target;
  assign icache_io_cpu_ras_update_bits_prediction_bits_entry = core_io_imem_ras_update_bits_prediction_bits_entry;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_history = core_io_imem_ras_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_value = core_io_imem_ras_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_flush_icache = core_io_imem_flush_icache;
  assign icache_io_cpu_flush_tlb = core_io_imem_flush_tlb;
  assign icache_io_ptw_req_ready = GEN_80;
  assign icache_io_ptw_resp_valid = GEN_81;
  assign icache_io_ptw_resp_bits_pte_reserved_for_hardware = GEN_82;
  assign icache_io_ptw_resp_bits_pte_ppn = GEN_83;
  assign icache_io_ptw_resp_bits_pte_reserved_for_software = GEN_84;
  assign icache_io_ptw_resp_bits_pte_d = GEN_85;
  assign icache_io_ptw_resp_bits_pte_a = GEN_86;
  assign icache_io_ptw_resp_bits_pte_g = GEN_87;
  assign icache_io_ptw_resp_bits_pte_u = GEN_88;
  assign icache_io_ptw_resp_bits_pte_x = GEN_89;
  assign icache_io_ptw_resp_bits_pte_w = GEN_90;
  assign icache_io_ptw_resp_bits_pte_r = GEN_91;
  assign icache_io_ptw_resp_bits_pte_v = GEN_92;
  assign icache_io_ptw_ptbr_asid = GEN_93;
  assign icache_io_ptw_ptbr_ppn = GEN_94;
  assign icache_io_ptw_invalidate = GEN_95;
  assign icache_io_ptw_status_debug = GEN_96;
  assign icache_io_ptw_status_prv = GEN_97;
  assign icache_io_ptw_status_sd = GEN_98;
  assign icache_io_ptw_status_zero3 = GEN_99;
  assign icache_io_ptw_status_sd_rv32 = GEN_100;
  assign icache_io_ptw_status_zero2 = GEN_101;
  assign icache_io_ptw_status_vm = GEN_102;
  assign icache_io_ptw_status_zero1 = GEN_103;
  assign icache_io_ptw_status_mxr = GEN_104;
  assign icache_io_ptw_status_pum = GEN_105;
  assign icache_io_ptw_status_mprv = GEN_106;
  assign icache_io_ptw_status_xs = GEN_107;
  assign icache_io_ptw_status_fs = GEN_108;
  assign icache_io_ptw_status_mpp = GEN_109;
  assign icache_io_ptw_status_hpp = GEN_110;
  assign icache_io_ptw_status_spp = GEN_111;
  assign icache_io_ptw_status_mpie = GEN_112;
  assign icache_io_ptw_status_hpie = GEN_113;
  assign icache_io_ptw_status_spie = GEN_114;
  assign icache_io_ptw_status_upie = GEN_115;
  assign icache_io_ptw_status_mie = GEN_116;
  assign icache_io_ptw_status_hie = GEN_117;
  assign icache_io_ptw_status_sie = GEN_118;
  assign icache_io_ptw_status_uie = GEN_119;
  assign icache_io_mem_acquire_ready = uncachedArb_io_in_0_acquire_ready;
  assign icache_io_mem_grant_valid = uncachedArb_io_in_0_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = uncachedArb_io_in_0_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = uncachedArb_io_in_0_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = uncachedArb_io_in_0_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = uncachedArb_io_in_0_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = uncachedArb_io_in_0_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = uncachedArb_io_in_0_grant_bits_data;
  assign DCache_1_clk = clk;
  assign DCache_1_reset = reset;
  assign DCache_1_io_cpu_req_valid = dcArb_io_mem_req_valid;
  assign DCache_1_io_cpu_req_bits_addr = dcArb_io_mem_req_bits_addr;
  assign DCache_1_io_cpu_req_bits_tag = dcArb_io_mem_req_bits_tag;
  assign DCache_1_io_cpu_req_bits_cmd = dcArb_io_mem_req_bits_cmd;
  assign DCache_1_io_cpu_req_bits_typ = dcArb_io_mem_req_bits_typ;
  assign DCache_1_io_cpu_req_bits_phys = dcArb_io_mem_req_bits_phys;
  assign DCache_1_io_cpu_req_bits_data = dcArb_io_mem_req_bits_data;
  assign DCache_1_io_cpu_s1_kill = dcArb_io_mem_s1_kill;
  assign DCache_1_io_cpu_s1_data = dcArb_io_mem_s1_data;
  assign DCache_1_io_cpu_invalidate_lr = dcArb_io_mem_invalidate_lr;
  assign DCache_1_io_ptw_req_ready = GEN_120;
  assign DCache_1_io_ptw_resp_valid = GEN_121;
  assign DCache_1_io_ptw_resp_bits_pte_reserved_for_hardware = GEN_122;
  assign DCache_1_io_ptw_resp_bits_pte_ppn = GEN_123;
  assign DCache_1_io_ptw_resp_bits_pte_reserved_for_software = GEN_124;
  assign DCache_1_io_ptw_resp_bits_pte_d = GEN_125;
  assign DCache_1_io_ptw_resp_bits_pte_a = GEN_126;
  assign DCache_1_io_ptw_resp_bits_pte_g = GEN_127;
  assign DCache_1_io_ptw_resp_bits_pte_u = GEN_128;
  assign DCache_1_io_ptw_resp_bits_pte_x = GEN_129;
  assign DCache_1_io_ptw_resp_bits_pte_w = GEN_130;
  assign DCache_1_io_ptw_resp_bits_pte_r = GEN_131;
  assign DCache_1_io_ptw_resp_bits_pte_v = GEN_132;
  assign DCache_1_io_ptw_ptbr_asid = GEN_133;
  assign DCache_1_io_ptw_ptbr_ppn = GEN_134;
  assign DCache_1_io_ptw_invalidate = GEN_135;
  assign DCache_1_io_ptw_status_debug = GEN_136;
  assign DCache_1_io_ptw_status_prv = GEN_137;
  assign DCache_1_io_ptw_status_sd = GEN_138;
  assign DCache_1_io_ptw_status_zero3 = GEN_139;
  assign DCache_1_io_ptw_status_sd_rv32 = GEN_140;
  assign DCache_1_io_ptw_status_zero2 = GEN_141;
  assign DCache_1_io_ptw_status_vm = GEN_142;
  assign DCache_1_io_ptw_status_zero1 = GEN_143;
  assign DCache_1_io_ptw_status_mxr = GEN_144;
  assign DCache_1_io_ptw_status_pum = GEN_145;
  assign DCache_1_io_ptw_status_mprv = GEN_146;
  assign DCache_1_io_ptw_status_xs = GEN_147;
  assign DCache_1_io_ptw_status_fs = GEN_148;
  assign DCache_1_io_ptw_status_mpp = GEN_149;
  assign DCache_1_io_ptw_status_hpp = GEN_150;
  assign DCache_1_io_ptw_status_spp = GEN_151;
  assign DCache_1_io_ptw_status_mpie = GEN_152;
  assign DCache_1_io_ptw_status_hpie = GEN_153;
  assign DCache_1_io_ptw_status_spie = GEN_154;
  assign DCache_1_io_ptw_status_upie = GEN_155;
  assign DCache_1_io_ptw_status_mie = GEN_156;
  assign DCache_1_io_ptw_status_hie = GEN_157;
  assign DCache_1_io_ptw_status_sie = GEN_158;
  assign DCache_1_io_ptw_status_uie = GEN_159;
  assign DCache_1_io_mem_acquire_ready = io_cached_0_acquire_ready;
  assign DCache_1_io_mem_probe_valid = io_cached_0_probe_valid;
  assign DCache_1_io_mem_probe_bits_addr_block = io_cached_0_probe_bits_addr_block;
  assign DCache_1_io_mem_probe_bits_p_type = io_cached_0_probe_bits_p_type;
  assign DCache_1_io_mem_release_ready = io_cached_0_release_ready;
  assign DCache_1_io_mem_grant_valid = io_cached_0_grant_valid;
  assign DCache_1_io_mem_grant_bits_addr_beat = io_cached_0_grant_bits_addr_beat;
  assign DCache_1_io_mem_grant_bits_client_xact_id = io_cached_0_grant_bits_client_xact_id;
  assign DCache_1_io_mem_grant_bits_manager_xact_id = io_cached_0_grant_bits_manager_xact_id;
  assign DCache_1_io_mem_grant_bits_is_builtin_type = io_cached_0_grant_bits_is_builtin_type;
  assign DCache_1_io_mem_grant_bits_g_type = io_cached_0_grant_bits_g_type;
  assign DCache_1_io_mem_grant_bits_data = io_cached_0_grant_bits_data;
  assign DCache_1_io_mem_grant_bits_manager_id = io_cached_0_grant_bits_manager_id;
  assign DCache_1_io_mem_finish_ready = io_cached_0_finish_ready;
  assign uncachedArb_clk = clk;
  assign uncachedArb_reset = reset;
  assign uncachedArb_io_in_0_acquire_valid = icache_io_mem_acquire_valid;
  assign uncachedArb_io_in_0_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign uncachedArb_io_in_0_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign uncachedArb_io_in_0_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign uncachedArb_io_in_0_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign uncachedArb_io_in_0_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign uncachedArb_io_in_0_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign uncachedArb_io_in_0_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign uncachedArb_io_in_0_grant_ready = icache_io_mem_grant_ready;
  assign uncachedArb_io_out_acquire_ready = io_uncached_0_acquire_ready;
  assign uncachedArb_io_out_grant_valid = io_uncached_0_grant_valid;
  assign uncachedArb_io_out_grant_bits_addr_beat = io_uncached_0_grant_bits_addr_beat;
  assign uncachedArb_io_out_grant_bits_client_xact_id = io_uncached_0_grant_bits_client_xact_id;
  assign uncachedArb_io_out_grant_bits_manager_xact_id = io_uncached_0_grant_bits_manager_xact_id;
  assign uncachedArb_io_out_grant_bits_is_builtin_type = io_uncached_0_grant_bits_is_builtin_type;
  assign uncachedArb_io_out_grant_bits_g_type = io_uncached_0_grant_bits_g_type;
  assign uncachedArb_io_out_grant_bits_data = io_uncached_0_grant_bits_data;
  assign dcArb_clk = clk;
  assign dcArb_reset = reset;
  assign dcArb_io_requestor_0_req_valid = core_io_dmem_req_valid;
  assign dcArb_io_requestor_0_req_bits_addr = core_io_dmem_req_bits_addr;
  assign dcArb_io_requestor_0_req_bits_tag = core_io_dmem_req_bits_tag;
  assign dcArb_io_requestor_0_req_bits_cmd = core_io_dmem_req_bits_cmd;
  assign dcArb_io_requestor_0_req_bits_typ = core_io_dmem_req_bits_typ;
  assign dcArb_io_requestor_0_req_bits_phys = core_io_dmem_req_bits_phys;
  assign dcArb_io_requestor_0_req_bits_data = core_io_dmem_req_bits_data;
  assign dcArb_io_requestor_0_s1_kill = core_io_dmem_s1_kill;
  assign dcArb_io_requestor_0_s1_data = core_io_dmem_s1_data;
  assign dcArb_io_requestor_0_invalidate_lr = core_io_dmem_invalidate_lr;
  assign dcArb_io_mem_req_ready = DCache_1_io_cpu_req_ready;
  assign dcArb_io_mem_s2_nack = DCache_1_io_cpu_s2_nack;
  assign dcArb_io_mem_resp_valid = DCache_1_io_cpu_resp_valid;
  assign dcArb_io_mem_resp_bits_addr = DCache_1_io_cpu_resp_bits_addr;
  assign dcArb_io_mem_resp_bits_tag = DCache_1_io_cpu_resp_bits_tag;
  assign dcArb_io_mem_resp_bits_cmd = DCache_1_io_cpu_resp_bits_cmd;
  assign dcArb_io_mem_resp_bits_typ = DCache_1_io_cpu_resp_bits_typ;
  assign dcArb_io_mem_resp_bits_data = DCache_1_io_cpu_resp_bits_data;
  assign dcArb_io_mem_resp_bits_replay = DCache_1_io_cpu_resp_bits_replay;
  assign dcArb_io_mem_resp_bits_has_data = DCache_1_io_cpu_resp_bits_has_data;
  assign dcArb_io_mem_resp_bits_data_word_bypass = DCache_1_io_cpu_resp_bits_data_word_bypass;
  assign dcArb_io_mem_resp_bits_store_data = DCache_1_io_cpu_resp_bits_store_data;
  assign dcArb_io_mem_replay_next = DCache_1_io_cpu_replay_next;
  assign dcArb_io_mem_xcpt_ma_ld = DCache_1_io_cpu_xcpt_ma_ld;
  assign dcArb_io_mem_xcpt_ma_st = DCache_1_io_cpu_xcpt_ma_st;
  assign dcArb_io_mem_xcpt_pf_ld = DCache_1_io_cpu_xcpt_pf_ld;
  assign dcArb_io_mem_xcpt_pf_st = DCache_1_io_cpu_xcpt_pf_st;
  assign dcArb_io_mem_ordered = DCache_1_io_cpu_ordered;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_0 = GEN_160[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_161[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_162[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_163[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_4 = GEN_164[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_5 = GEN_165[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_6 = GEN_166[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_7 = GEN_167[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_8 = GEN_168[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_9 = GEN_169[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_10 = GEN_170[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_11 = GEN_171[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_12 = GEN_172[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_13 = GEN_173[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_14 = GEN_174[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_15 = GEN_175[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_16 = GEN_176[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_17 = GEN_177[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_18 = GEN_178[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_19 = GEN_179[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_20 = GEN_180[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_21 = GEN_181[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_22 = GEN_182[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_23 = GEN_183[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_24 = GEN_184[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_25 = GEN_185[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_26 = GEN_186[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_27 = GEN_187[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_28 = GEN_188[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_29 = GEN_189[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_190[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_191[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_32 = GEN_192[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_33 = GEN_193[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_34 = GEN_194[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_35 = GEN_195[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_36 = GEN_196[39:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_37 = GEN_197[5:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_38 = GEN_198[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_39 = GEN_199[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_40 = GEN_200[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_41 = GEN_201[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_42 = GEN_202[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_43 = GEN_203[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_44 = GEN_204[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_45 = GEN_205[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_46 = GEN_206[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_47 = GEN_207[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_48 = GEN_208[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_49 = GEN_209[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_50 = GEN_210[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_51 = GEN_211[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_52 = GEN_212[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_53 = GEN_213[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_54 = GEN_214[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_55 = GEN_215[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_56 = GEN_216[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_57 = GEN_217[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_58 = GEN_218[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_59 = GEN_219[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_60 = GEN_220[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_61 = GEN_221[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_62 = GEN_222[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_63 = GEN_223[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_64 = GEN_224[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_65 = GEN_225[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_66 = GEN_226[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_67 = GEN_227[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_68 = GEN_228[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_69 = GEN_229[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_70 = GEN_230[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_71 = GEN_231[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_72 = GEN_232[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_73 = GEN_233[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_74 = GEN_234[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_75 = GEN_235[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_76 = GEN_236[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_77 = GEN_237[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_78 = GEN_238[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_79 = GEN_239[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_80 = GEN_240[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_81 = GEN_241[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_82 = GEN_242[15:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_83 = GEN_243[37:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_84 = GEN_244[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_85 = GEN_245[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_86 = GEN_246[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_87 = GEN_247[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_88 = GEN_248[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_89 = GEN_249[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_90 = GEN_250[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_91 = GEN_251[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_92 = GEN_252[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_93 = GEN_253[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_94 = GEN_254[37:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_95 = GEN_255[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_96 = GEN_256[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_97 = GEN_257[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_98 = GEN_258[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_99 = GEN_259[30:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_100 = GEN_260[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_101 = GEN_261[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_102 = GEN_262[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_103 = GEN_263[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_104 = GEN_264[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_105 = GEN_265[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_106 = GEN_266[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_107 = GEN_267[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_108 = GEN_268[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_109 = GEN_269[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_110 = GEN_270[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_111 = GEN_271[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_112 = GEN_272[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_113 = GEN_273[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_114 = GEN_274[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_115 = GEN_275[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_116 = GEN_276[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_117 = GEN_277[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_118 = GEN_278[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_119 = GEN_279[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_120 = GEN_280[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_121 = GEN_281[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_122 = GEN_282[15:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_123 = GEN_283[37:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_124 = GEN_284[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_125 = GEN_285[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_126 = GEN_286[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_127 = GEN_287[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_128 = GEN_288[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_129 = GEN_289[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_130 = GEN_290[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_131 = GEN_291[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_132 = GEN_292[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_133 = GEN_293[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_134 = GEN_294[37:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_135 = GEN_295[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_136 = GEN_296[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_137 = GEN_297[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_138 = GEN_298[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_139 = GEN_299[30:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_140 = GEN_300[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_141 = GEN_301[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_142 = GEN_302[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_143 = GEN_303[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_144 = GEN_304[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_145 = GEN_305[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_146 = GEN_306[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_147 = GEN_307[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_148 = GEN_308[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_149 = GEN_309[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_150 = GEN_310[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_151 = GEN_311[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_152 = GEN_312[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_153 = GEN_313[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_154 = GEN_314[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_155 = GEN_315[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_156 = GEN_316[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_157 = GEN_317[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_158 = GEN_318[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_159 = GEN_319[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_160 = {1{$random}};
  GEN_161 = {1{$random}};
  GEN_162 = {2{$random}};
  GEN_163 = {2{$random}};
  GEN_164 = {1{$random}};
  GEN_165 = {1{$random}};
  GEN_166 = {1{$random}};
  GEN_167 = {1{$random}};
  GEN_168 = {1{$random}};
  GEN_169 = {1{$random}};
  GEN_170 = {1{$random}};
  GEN_171 = {1{$random}};
  GEN_172 = {1{$random}};
  GEN_173 = {1{$random}};
  GEN_174 = {1{$random}};
  GEN_175 = {1{$random}};
  GEN_176 = {1{$random}};
  GEN_177 = {1{$random}};
  GEN_178 = {1{$random}};
  GEN_179 = {1{$random}};
  GEN_180 = {1{$random}};
  GEN_181 = {1{$random}};
  GEN_182 = {1{$random}};
  GEN_183 = {1{$random}};
  GEN_184 = {1{$random}};
  GEN_185 = {1{$random}};
  GEN_186 = {1{$random}};
  GEN_187 = {1{$random}};
  GEN_188 = {1{$random}};
  GEN_189 = {3{$random}};
  GEN_190 = {1{$random}};
  GEN_191 = {1{$random}};
  GEN_192 = {1{$random}};
  GEN_193 = {1{$random}};
  GEN_194 = {2{$random}};
  GEN_195 = {1{$random}};
  GEN_196 = {2{$random}};
  GEN_197 = {1{$random}};
  GEN_198 = {1{$random}};
  GEN_199 = {1{$random}};
  GEN_200 = {1{$random}};
  GEN_201 = {2{$random}};
  GEN_202 = {1{$random}};
  GEN_203 = {2{$random}};
  GEN_204 = {1{$random}};
  GEN_205 = {1{$random}};
  GEN_206 = {1{$random}};
  GEN_207 = {1{$random}};
  GEN_208 = {1{$random}};
  GEN_209 = {1{$random}};
  GEN_210 = {1{$random}};
  GEN_211 = {1{$random}};
  GEN_212 = {1{$random}};
  GEN_213 = {1{$random}};
  GEN_214 = {2{$random}};
  GEN_215 = {1{$random}};
  GEN_216 = {1{$random}};
  GEN_217 = {1{$random}};
  GEN_218 = {1{$random}};
  GEN_219 = {1{$random}};
  GEN_220 = {1{$random}};
  GEN_221 = {1{$random}};
  GEN_222 = {1{$random}};
  GEN_223 = {1{$random}};
  GEN_224 = {1{$random}};
  GEN_225 = {1{$random}};
  GEN_226 = {1{$random}};
  GEN_227 = {1{$random}};
  GEN_228 = {1{$random}};
  GEN_229 = {1{$random}};
  GEN_230 = {1{$random}};
  GEN_231 = {1{$random}};
  GEN_232 = {1{$random}};
  GEN_233 = {1{$random}};
  GEN_234 = {1{$random}};
  GEN_235 = {1{$random}};
  GEN_236 = {3{$random}};
  GEN_237 = {3{$random}};
  GEN_238 = {3{$random}};
  GEN_239 = {1{$random}};
  GEN_240 = {1{$random}};
  GEN_241 = {1{$random}};
  GEN_242 = {1{$random}};
  GEN_243 = {2{$random}};
  GEN_244 = {1{$random}};
  GEN_245 = {1{$random}};
  GEN_246 = {1{$random}};
  GEN_247 = {1{$random}};
  GEN_248 = {1{$random}};
  GEN_249 = {1{$random}};
  GEN_250 = {1{$random}};
  GEN_251 = {1{$random}};
  GEN_252 = {1{$random}};
  GEN_253 = {1{$random}};
  GEN_254 = {2{$random}};
  GEN_255 = {1{$random}};
  GEN_256 = {1{$random}};
  GEN_257 = {1{$random}};
  GEN_258 = {1{$random}};
  GEN_259 = {1{$random}};
  GEN_260 = {1{$random}};
  GEN_261 = {1{$random}};
  GEN_262 = {1{$random}};
  GEN_263 = {1{$random}};
  GEN_264 = {1{$random}};
  GEN_265 = {1{$random}};
  GEN_266 = {1{$random}};
  GEN_267 = {1{$random}};
  GEN_268 = {1{$random}};
  GEN_269 = {1{$random}};
  GEN_270 = {1{$random}};
  GEN_271 = {1{$random}};
  GEN_272 = {1{$random}};
  GEN_273 = {1{$random}};
  GEN_274 = {1{$random}};
  GEN_275 = {1{$random}};
  GEN_276 = {1{$random}};
  GEN_277 = {1{$random}};
  GEN_278 = {1{$random}};
  GEN_279 = {1{$random}};
  GEN_280 = {1{$random}};
  GEN_281 = {1{$random}};
  GEN_282 = {1{$random}};
  GEN_283 = {2{$random}};
  GEN_284 = {1{$random}};
  GEN_285 = {1{$random}};
  GEN_286 = {1{$random}};
  GEN_287 = {1{$random}};
  GEN_288 = {1{$random}};
  GEN_289 = {1{$random}};
  GEN_290 = {1{$random}};
  GEN_291 = {1{$random}};
  GEN_292 = {1{$random}};
  GEN_293 = {1{$random}};
  GEN_294 = {2{$random}};
  GEN_295 = {1{$random}};
  GEN_296 = {1{$random}};
  GEN_297 = {1{$random}};
  GEN_298 = {1{$random}};
  GEN_299 = {1{$random}};
  GEN_300 = {1{$random}};
  GEN_301 = {1{$random}};
  GEN_302 = {1{$random}};
  GEN_303 = {1{$random}};
  GEN_304 = {1{$random}};
  GEN_305 = {1{$random}};
  GEN_306 = {1{$random}};
  GEN_307 = {1{$random}};
  GEN_308 = {1{$random}};
  GEN_309 = {1{$random}};
  GEN_310 = {1{$random}};
  GEN_311 = {1{$random}};
  GEN_312 = {1{$random}};
  GEN_313 = {1{$random}};
  GEN_314 = {1{$random}};
  GEN_315 = {1{$random}};
  GEN_316 = {1{$random}};
  GEN_317 = {1{$random}};
  GEN_318 = {1{$random}};
  GEN_319 = {1{$random}};
  end
`endif
endmodule
module Queue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input   io_enq_bits_payload_client_xact_id,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input   io_enq_bits_payload_is_builtin_type,
  input  [2:0] io_enq_bits_payload_a_type,
  input  [10:0] io_enq_bits_payload_union,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output  io_deq_bits_payload_client_xact_id,
  output [2:0] io_deq_bits_payload_addr_beat,
  output  io_deq_bits_payload_is_builtin_type,
  output [2:0] io_deq_bits_payload_a_type,
  output [10:0] io_deq_bits_payload_union,
  output [63:0] io_deq_bits_payload_data,
  output  io_count
);
  reg [1:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1144_data;
  wire  ram_header_src_T_1144_addr;
  wire  ram_header_src_T_1144_en;
  wire [1:0] ram_header_src_T_1025_data;
  wire  ram_header_src_T_1025_addr;
  wire  ram_header_src_T_1025_mask;
  wire  ram_header_src_T_1025_en;
  reg [1:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1144_data;
  wire  ram_header_dst_T_1144_addr;
  wire  ram_header_dst_T_1144_en;
  wire [1:0] ram_header_dst_T_1025_data;
  wire  ram_header_dst_T_1025_addr;
  wire  ram_header_dst_T_1025_mask;
  wire  ram_header_dst_T_1025_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1144_data;
  wire  ram_payload_addr_block_T_1144_addr;
  wire  ram_payload_addr_block_T_1144_en;
  wire [25:0] ram_payload_addr_block_T_1025_data;
  wire  ram_payload_addr_block_T_1025_addr;
  wire  ram_payload_addr_block_T_1025_mask;
  wire  ram_payload_addr_block_T_1025_en;
  reg  ram_payload_client_xact_id [0:0];
  reg [31:0] GEN_3;
  wire  ram_payload_client_xact_id_T_1144_data;
  wire  ram_payload_client_xact_id_T_1144_addr;
  wire  ram_payload_client_xact_id_T_1144_en;
  wire  ram_payload_client_xact_id_T_1025_data;
  wire  ram_payload_client_xact_id_T_1025_addr;
  wire  ram_payload_client_xact_id_T_1025_mask;
  wire  ram_payload_client_xact_id_T_1025_en;
  reg [2:0] ram_payload_addr_beat [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_payload_addr_beat_T_1144_data;
  wire  ram_payload_addr_beat_T_1144_addr;
  wire  ram_payload_addr_beat_T_1144_en;
  wire [2:0] ram_payload_addr_beat_T_1025_data;
  wire  ram_payload_addr_beat_T_1025_addr;
  wire  ram_payload_addr_beat_T_1025_mask;
  wire  ram_payload_addr_beat_T_1025_en;
  reg  ram_payload_is_builtin_type [0:0];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1144_data;
  wire  ram_payload_is_builtin_type_T_1144_addr;
  wire  ram_payload_is_builtin_type_T_1144_en;
  wire  ram_payload_is_builtin_type_T_1025_data;
  wire  ram_payload_is_builtin_type_T_1025_addr;
  wire  ram_payload_is_builtin_type_T_1025_mask;
  wire  ram_payload_is_builtin_type_T_1025_en;
  reg [2:0] ram_payload_a_type [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_a_type_T_1144_data;
  wire  ram_payload_a_type_T_1144_addr;
  wire  ram_payload_a_type_T_1144_en;
  wire [2:0] ram_payload_a_type_T_1025_data;
  wire  ram_payload_a_type_T_1025_addr;
  wire  ram_payload_a_type_T_1025_mask;
  wire  ram_payload_a_type_T_1025_en;
  reg [10:0] ram_payload_union [0:0];
  reg [31:0] GEN_7;
  wire [10:0] ram_payload_union_T_1144_data;
  wire  ram_payload_union_T_1144_addr;
  wire  ram_payload_union_T_1144_en;
  wire [10:0] ram_payload_union_T_1025_data;
  wire  ram_payload_union_T_1025_addr;
  wire  ram_payload_union_T_1025_mask;
  wire  ram_payload_union_T_1025_en;
  reg [63:0] ram_payload_data [0:0];
  reg [63:0] GEN_8;
  wire [63:0] ram_payload_data_T_1144_data;
  wire  ram_payload_data_T_1144_addr;
  wire  ram_payload_data_T_1144_en;
  wire [63:0] ram_payload_data_T_1025_data;
  wire  ram_payload_data_T_1025_addr;
  wire  ram_payload_data_T_1025_mask;
  wire  ram_payload_data_T_1025_en;
  reg  maybe_full;
  reg [31:0] GEN_9;
  wire  T_1022;
  wire  T_1023;
  wire  do_enq;
  wire  T_1024;
  wire  do_deq;
  wire  T_1139;
  wire  GEN_21;
  wire  T_1141;
  wire [1:0] T_1256;
  wire  ptr_diff;
  wire [1:0] T_1258;
  assign io_enq_ready = T_1022;
  assign io_deq_valid = T_1141;
  assign io_deq_bits_header_src = ram_header_src_T_1144_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1144_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1144_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1144_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1144_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1144_data;
  assign io_deq_bits_payload_a_type = ram_payload_a_type_T_1144_data;
  assign io_deq_bits_payload_union = ram_payload_union_T_1144_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1144_data;
  assign io_count = T_1258[0];
  assign ram_header_src_T_1144_addr = 1'h0;
  assign ram_header_src_T_1144_en = 1'h1;
  assign ram_header_src_T_1144_data = ram_header_src[ram_header_src_T_1144_addr];
  assign ram_header_src_T_1025_data = io_enq_bits_header_src;
  assign ram_header_src_T_1025_addr = 1'h0;
  assign ram_header_src_T_1025_mask = do_enq;
  assign ram_header_src_T_1025_en = do_enq;
  assign ram_header_dst_T_1144_addr = 1'h0;
  assign ram_header_dst_T_1144_en = 1'h1;
  assign ram_header_dst_T_1144_data = ram_header_dst[ram_header_dst_T_1144_addr];
  assign ram_header_dst_T_1025_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1025_addr = 1'h0;
  assign ram_header_dst_T_1025_mask = do_enq;
  assign ram_header_dst_T_1025_en = do_enq;
  assign ram_payload_addr_block_T_1144_addr = 1'h0;
  assign ram_payload_addr_block_T_1144_en = 1'h1;
  assign ram_payload_addr_block_T_1144_data = ram_payload_addr_block[ram_payload_addr_block_T_1144_addr];
  assign ram_payload_addr_block_T_1025_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1025_addr = 1'h0;
  assign ram_payload_addr_block_T_1025_mask = do_enq;
  assign ram_payload_addr_block_T_1025_en = do_enq;
  assign ram_payload_client_xact_id_T_1144_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1144_en = 1'h1;
  assign ram_payload_client_xact_id_T_1144_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1144_addr];
  assign ram_payload_client_xact_id_T_1025_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1025_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1025_mask = do_enq;
  assign ram_payload_client_xact_id_T_1025_en = do_enq;
  assign ram_payload_addr_beat_T_1144_addr = 1'h0;
  assign ram_payload_addr_beat_T_1144_en = 1'h1;
  assign ram_payload_addr_beat_T_1144_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1144_addr];
  assign ram_payload_addr_beat_T_1025_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1025_addr = 1'h0;
  assign ram_payload_addr_beat_T_1025_mask = do_enq;
  assign ram_payload_addr_beat_T_1025_en = do_enq;
  assign ram_payload_is_builtin_type_T_1144_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1144_en = 1'h1;
  assign ram_payload_is_builtin_type_T_1144_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1144_addr];
  assign ram_payload_is_builtin_type_T_1025_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1025_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1025_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1025_en = do_enq;
  assign ram_payload_a_type_T_1144_addr = 1'h0;
  assign ram_payload_a_type_T_1144_en = 1'h1;
  assign ram_payload_a_type_T_1144_data = ram_payload_a_type[ram_payload_a_type_T_1144_addr];
  assign ram_payload_a_type_T_1025_data = io_enq_bits_payload_a_type;
  assign ram_payload_a_type_T_1025_addr = 1'h0;
  assign ram_payload_a_type_T_1025_mask = do_enq;
  assign ram_payload_a_type_T_1025_en = do_enq;
  assign ram_payload_union_T_1144_addr = 1'h0;
  assign ram_payload_union_T_1144_en = 1'h1;
  assign ram_payload_union_T_1144_data = ram_payload_union[ram_payload_union_T_1144_addr];
  assign ram_payload_union_T_1025_data = io_enq_bits_payload_union;
  assign ram_payload_union_T_1025_addr = 1'h0;
  assign ram_payload_union_T_1025_mask = do_enq;
  assign ram_payload_union_T_1025_en = do_enq;
  assign ram_payload_data_T_1144_addr = 1'h0;
  assign ram_payload_data_T_1144_en = 1'h1;
  assign ram_payload_data_T_1144_data = ram_payload_data[ram_payload_data_T_1144_addr];
  assign ram_payload_data_T_1025_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1025_addr = 1'h0;
  assign ram_payload_data_T_1025_mask = do_enq;
  assign ram_payload_data_T_1025_en = do_enq;
  assign T_1022 = maybe_full == 1'h0;
  assign T_1023 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1023;
  assign T_1024 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1024;
  assign T_1139 = do_enq != do_deq;
  assign GEN_21 = T_1139 ? do_enq : maybe_full;
  assign T_1141 = T_1022 == 1'h0;
  assign T_1256 = 1'h0 - 1'h0;
  assign ptr_diff = T_1256[0:0];
  assign T_1258 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_4[2:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_a_type[initvar] = GEN_6[2:0];
  `endif
  GEN_7 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_union[initvar] = GEN_7[10:0];
  `endif
  GEN_8 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_8[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {1{$random}};
  maybe_full = GEN_9[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1025_en & ram_header_src_T_1025_mask) begin
      ram_header_src[ram_header_src_T_1025_addr] <= ram_header_src_T_1025_data;
    end
    if(ram_header_dst_T_1025_en & ram_header_dst_T_1025_mask) begin
      ram_header_dst[ram_header_dst_T_1025_addr] <= ram_header_dst_T_1025_data;
    end
    if(ram_payload_addr_block_T_1025_en & ram_payload_addr_block_T_1025_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1025_addr] <= ram_payload_addr_block_T_1025_data;
    end
    if(ram_payload_client_xact_id_T_1025_en & ram_payload_client_xact_id_T_1025_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1025_addr] <= ram_payload_client_xact_id_T_1025_data;
    end
    if(ram_payload_addr_beat_T_1025_en & ram_payload_addr_beat_T_1025_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1025_addr] <= ram_payload_addr_beat_T_1025_data;
    end
    if(ram_payload_is_builtin_type_T_1025_en & ram_payload_is_builtin_type_T_1025_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1025_addr] <= ram_payload_is_builtin_type_T_1025_data;
    end
    if(ram_payload_a_type_T_1025_en & ram_payload_a_type_T_1025_mask) begin
      ram_payload_a_type[ram_payload_a_type_T_1025_addr] <= ram_payload_a_type_T_1025_data;
    end
    if(ram_payload_union_T_1025_en & ram_payload_union_T_1025_mask) begin
      ram_payload_union[ram_payload_union_T_1025_addr] <= ram_payload_union_T_1025_data;
    end
    if(ram_payload_data_T_1025_en & ram_payload_data_T_1025_mask) begin
      ram_payload_data[ram_payload_data_T_1025_addr] <= ram_payload_data_T_1025_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_1(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_p_type,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_p_type,
  output  io_count
);
  reg [1:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1094_data;
  wire  ram_header_src_T_1094_addr;
  wire  ram_header_src_T_1094_en;
  wire [1:0] ram_header_src_T_980_data;
  wire  ram_header_src_T_980_addr;
  wire  ram_header_src_T_980_mask;
  wire  ram_header_src_T_980_en;
  reg [1:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1094_data;
  wire  ram_header_dst_T_1094_addr;
  wire  ram_header_dst_T_1094_en;
  wire [1:0] ram_header_dst_T_980_data;
  wire  ram_header_dst_T_980_addr;
  wire  ram_header_dst_T_980_mask;
  wire  ram_header_dst_T_980_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1094_data;
  wire  ram_payload_addr_block_T_1094_addr;
  wire  ram_payload_addr_block_T_1094_en;
  wire [25:0] ram_payload_addr_block_T_980_data;
  wire  ram_payload_addr_block_T_980_addr;
  wire  ram_payload_addr_block_T_980_mask;
  wire  ram_payload_addr_block_T_980_en;
  reg [1:0] ram_payload_p_type [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_p_type_T_1094_data;
  wire  ram_payload_p_type_T_1094_addr;
  wire  ram_payload_p_type_T_1094_en;
  wire [1:0] ram_payload_p_type_T_980_data;
  wire  ram_payload_p_type_T_980_addr;
  wire  ram_payload_p_type_T_980_mask;
  wire  ram_payload_p_type_T_980_en;
  reg  maybe_full;
  reg [31:0] GEN_4;
  wire  T_977;
  wire  T_978;
  wire  do_enq;
  wire  T_979;
  wire  do_deq;
  wire  T_1089;
  wire  GEN_11;
  wire  T_1091;
  wire [1:0] T_1201;
  wire  ptr_diff;
  wire [1:0] T_1203;
  assign io_enq_ready = T_977;
  assign io_deq_valid = T_1091;
  assign io_deq_bits_header_src = ram_header_src_T_1094_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1094_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1094_data;
  assign io_deq_bits_payload_p_type = ram_payload_p_type_T_1094_data;
  assign io_count = T_1203[0];
  assign ram_header_src_T_1094_addr = 1'h0;
  assign ram_header_src_T_1094_en = 1'h1;
  assign ram_header_src_T_1094_data = ram_header_src[ram_header_src_T_1094_addr];
  assign ram_header_src_T_980_data = io_enq_bits_header_src;
  assign ram_header_src_T_980_addr = 1'h0;
  assign ram_header_src_T_980_mask = do_enq;
  assign ram_header_src_T_980_en = do_enq;
  assign ram_header_dst_T_1094_addr = 1'h0;
  assign ram_header_dst_T_1094_en = 1'h1;
  assign ram_header_dst_T_1094_data = ram_header_dst[ram_header_dst_T_1094_addr];
  assign ram_header_dst_T_980_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_980_addr = 1'h0;
  assign ram_header_dst_T_980_mask = do_enq;
  assign ram_header_dst_T_980_en = do_enq;
  assign ram_payload_addr_block_T_1094_addr = 1'h0;
  assign ram_payload_addr_block_T_1094_en = 1'h1;
  assign ram_payload_addr_block_T_1094_data = ram_payload_addr_block[ram_payload_addr_block_T_1094_addr];
  assign ram_payload_addr_block_T_980_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_980_addr = 1'h0;
  assign ram_payload_addr_block_T_980_mask = do_enq;
  assign ram_payload_addr_block_T_980_en = do_enq;
  assign ram_payload_p_type_T_1094_addr = 1'h0;
  assign ram_payload_p_type_T_1094_en = 1'h1;
  assign ram_payload_p_type_T_1094_data = ram_payload_p_type[ram_payload_p_type_T_1094_addr];
  assign ram_payload_p_type_T_980_data = io_enq_bits_payload_p_type;
  assign ram_payload_p_type_T_980_addr = 1'h0;
  assign ram_payload_p_type_T_980_mask = do_enq;
  assign ram_payload_p_type_T_980_en = do_enq;
  assign T_977 = maybe_full == 1'h0;
  assign T_978 = io_enq_ready & io_enq_valid;
  assign do_enq = T_978;
  assign T_979 = io_deq_ready & io_deq_valid;
  assign do_deq = T_979;
  assign T_1089 = do_enq != do_deq;
  assign GEN_11 = T_1089 ? do_enq : maybe_full;
  assign T_1091 = T_977 == 1'h0;
  assign T_1201 = 1'h0 - 1'h0;
  assign ptr_diff = T_1201[0:0];
  assign T_1203 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_p_type[initvar] = GEN_3[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {1{$random}};
  maybe_full = GEN_4[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_980_en & ram_header_src_T_980_mask) begin
      ram_header_src[ram_header_src_T_980_addr] <= ram_header_src_T_980_data;
    end
    if(ram_header_dst_T_980_en & ram_header_dst_T_980_mask) begin
      ram_header_dst[ram_header_dst_T_980_addr] <= ram_header_dst_T_980_data;
    end
    if(ram_payload_addr_block_T_980_en & ram_payload_addr_block_T_980_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_980_addr] <= ram_payload_addr_block_T_980_data;
    end
    if(ram_payload_p_type_T_980_en & ram_payload_p_type_T_980_mask) begin
      ram_payload_p_type[ram_payload_p_type_T_980_addr] <= ram_payload_p_type_T_980_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1089) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_2(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input  [25:0] io_enq_bits_payload_addr_block,
  input   io_enq_bits_payload_client_xact_id,
  input   io_enq_bits_payload_voluntary,
  input  [2:0] io_enq_bits_payload_r_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output [25:0] io_deq_bits_payload_addr_block,
  output  io_deq_bits_payload_client_xact_id,
  output  io_deq_bits_payload_voluntary,
  output [2:0] io_deq_bits_payload_r_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [1:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1144_data;
  wire  ram_header_src_T_1144_addr;
  wire  ram_header_src_T_1144_en;
  wire [1:0] ram_header_src_T_1018_data;
  wire  ram_header_src_T_1018_addr;
  wire  ram_header_src_T_1018_mask;
  wire  ram_header_src_T_1018_en;
  reg [1:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1144_data;
  wire  ram_header_dst_T_1144_addr;
  wire  ram_header_dst_T_1144_en;
  wire [1:0] ram_header_dst_T_1018_data;
  wire  ram_header_dst_T_1018_addr;
  wire  ram_header_dst_T_1018_mask;
  wire  ram_header_dst_T_1018_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1144_data;
  wire  ram_payload_addr_beat_T_1144_addr;
  wire  ram_payload_addr_beat_T_1144_en;
  wire [2:0] ram_payload_addr_beat_T_1018_data;
  wire  ram_payload_addr_beat_T_1018_addr;
  wire  ram_payload_addr_beat_T_1018_mask;
  wire  ram_payload_addr_beat_T_1018_en;
  reg [25:0] ram_payload_addr_block [0:1];
  reg [31:0] GEN_3;
  wire [25:0] ram_payload_addr_block_T_1144_data;
  wire  ram_payload_addr_block_T_1144_addr;
  wire  ram_payload_addr_block_T_1144_en;
  wire [25:0] ram_payload_addr_block_T_1018_data;
  wire  ram_payload_addr_block_T_1018_addr;
  wire  ram_payload_addr_block_T_1018_mask;
  wire  ram_payload_addr_block_T_1018_en;
  reg  ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_4;
  wire  ram_payload_client_xact_id_T_1144_data;
  wire  ram_payload_client_xact_id_T_1144_addr;
  wire  ram_payload_client_xact_id_T_1144_en;
  wire  ram_payload_client_xact_id_T_1018_data;
  wire  ram_payload_client_xact_id_T_1018_addr;
  wire  ram_payload_client_xact_id_T_1018_mask;
  wire  ram_payload_client_xact_id_T_1018_en;
  reg  ram_payload_voluntary [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_voluntary_T_1144_data;
  wire  ram_payload_voluntary_T_1144_addr;
  wire  ram_payload_voluntary_T_1144_en;
  wire  ram_payload_voluntary_T_1018_data;
  wire  ram_payload_voluntary_T_1018_addr;
  wire  ram_payload_voluntary_T_1018_mask;
  wire  ram_payload_voluntary_T_1018_en;
  reg [2:0] ram_payload_r_type [0:1];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_r_type_T_1144_data;
  wire  ram_payload_r_type_T_1144_addr;
  wire  ram_payload_r_type_T_1144_en;
  wire [2:0] ram_payload_r_type_T_1018_data;
  wire  ram_payload_r_type_T_1018_addr;
  wire  ram_payload_r_type_T_1018_mask;
  wire  ram_payload_r_type_T_1018_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1144_data;
  wire  ram_payload_data_T_1144_addr;
  wire  ram_payload_data_T_1144_en;
  wire [63:0] ram_payload_data_T_1018_data;
  wire  ram_payload_data_T_1018_addr;
  wire  ram_payload_data_T_1018_mask;
  wire  ram_payload_data_T_1018_en;
  reg  T_1010;
  reg [31:0] GEN_8;
  reg  T_1012;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1015;
  wire  empty;
  wire  full;
  wire  T_1016;
  wire  do_enq;
  wire  T_1017;
  wire  do_deq;
  wire [1:0] T_1132;
  wire  T_1133;
  wire  GEN_19;
  wire [1:0] T_1137;
  wire  T_1138;
  wire  GEN_20;
  wire  T_1139;
  wire  GEN_21;
  wire  T_1141;
  wire  T_1143;
  wire [1:0] T_1255;
  wire  ptr_diff;
  wire  T_1256;
  wire [1:0] T_1257;
  assign io_enq_ready = T_1143;
  assign io_deq_valid = T_1141;
  assign io_deq_bits_header_src = ram_header_src_T_1144_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1144_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1144_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1144_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1144_data;
  assign io_deq_bits_payload_voluntary = ram_payload_voluntary_T_1144_data;
  assign io_deq_bits_payload_r_type = ram_payload_r_type_T_1144_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1144_data;
  assign io_count = T_1257;
  assign ram_header_src_T_1144_addr = T_1012;
  assign ram_header_src_T_1144_en = 1'h1;
  assign ram_header_src_T_1144_data = ram_header_src[ram_header_src_T_1144_addr];
  assign ram_header_src_T_1018_data = io_enq_bits_header_src;
  assign ram_header_src_T_1018_addr = T_1010;
  assign ram_header_src_T_1018_mask = do_enq;
  assign ram_header_src_T_1018_en = do_enq;
  assign ram_header_dst_T_1144_addr = T_1012;
  assign ram_header_dst_T_1144_en = 1'h1;
  assign ram_header_dst_T_1144_data = ram_header_dst[ram_header_dst_T_1144_addr];
  assign ram_header_dst_T_1018_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1018_addr = T_1010;
  assign ram_header_dst_T_1018_mask = do_enq;
  assign ram_header_dst_T_1018_en = do_enq;
  assign ram_payload_addr_beat_T_1144_addr = T_1012;
  assign ram_payload_addr_beat_T_1144_en = 1'h1;
  assign ram_payload_addr_beat_T_1144_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1144_addr];
  assign ram_payload_addr_beat_T_1018_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1018_addr = T_1010;
  assign ram_payload_addr_beat_T_1018_mask = do_enq;
  assign ram_payload_addr_beat_T_1018_en = do_enq;
  assign ram_payload_addr_block_T_1144_addr = T_1012;
  assign ram_payload_addr_block_T_1144_en = 1'h1;
  assign ram_payload_addr_block_T_1144_data = ram_payload_addr_block[ram_payload_addr_block_T_1144_addr];
  assign ram_payload_addr_block_T_1018_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1018_addr = T_1010;
  assign ram_payload_addr_block_T_1018_mask = do_enq;
  assign ram_payload_addr_block_T_1018_en = do_enq;
  assign ram_payload_client_xact_id_T_1144_addr = T_1012;
  assign ram_payload_client_xact_id_T_1144_en = 1'h1;
  assign ram_payload_client_xact_id_T_1144_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1144_addr];
  assign ram_payload_client_xact_id_T_1018_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1018_addr = T_1010;
  assign ram_payload_client_xact_id_T_1018_mask = do_enq;
  assign ram_payload_client_xact_id_T_1018_en = do_enq;
  assign ram_payload_voluntary_T_1144_addr = T_1012;
  assign ram_payload_voluntary_T_1144_en = 1'h1;
  assign ram_payload_voluntary_T_1144_data = ram_payload_voluntary[ram_payload_voluntary_T_1144_addr];
  assign ram_payload_voluntary_T_1018_data = io_enq_bits_payload_voluntary;
  assign ram_payload_voluntary_T_1018_addr = T_1010;
  assign ram_payload_voluntary_T_1018_mask = do_enq;
  assign ram_payload_voluntary_T_1018_en = do_enq;
  assign ram_payload_r_type_T_1144_addr = T_1012;
  assign ram_payload_r_type_T_1144_en = 1'h1;
  assign ram_payload_r_type_T_1144_data = ram_payload_r_type[ram_payload_r_type_T_1144_addr];
  assign ram_payload_r_type_T_1018_data = io_enq_bits_payload_r_type;
  assign ram_payload_r_type_T_1018_addr = T_1010;
  assign ram_payload_r_type_T_1018_mask = do_enq;
  assign ram_payload_r_type_T_1018_en = do_enq;
  assign ram_payload_data_T_1144_addr = T_1012;
  assign ram_payload_data_T_1144_en = 1'h1;
  assign ram_payload_data_T_1144_data = ram_payload_data[ram_payload_data_T_1144_addr];
  assign ram_payload_data_T_1018_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1018_addr = T_1010;
  assign ram_payload_data_T_1018_mask = do_enq;
  assign ram_payload_data_T_1018_en = do_enq;
  assign ptr_match = T_1010 == T_1012;
  assign T_1015 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1015;
  assign full = ptr_match & maybe_full;
  assign T_1016 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1016;
  assign T_1017 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1017;
  assign T_1132 = T_1010 + 1'h1;
  assign T_1133 = T_1132[0:0];
  assign GEN_19 = do_enq ? T_1133 : T_1010;
  assign T_1137 = T_1012 + 1'h1;
  assign T_1138 = T_1137[0:0];
  assign GEN_20 = do_deq ? T_1138 : T_1012;
  assign T_1139 = do_enq != do_deq;
  assign GEN_21 = T_1139 ? do_enq : maybe_full;
  assign T_1141 = empty == 1'h0;
  assign T_1143 = full == 1'h0;
  assign T_1255 = T_1010 - T_1012;
  assign ptr_diff = T_1255[0:0];
  assign T_1256 = maybe_full & ptr_match;
  assign T_1257 = {T_1256,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_3[25:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_4[0:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_voluntary[initvar] = GEN_5[0:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_r_type[initvar] = GEN_6[2:0];
  `endif
  GEN_7 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  T_1010 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {1{$random}};
  T_1012 = GEN_9[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1018_en & ram_header_src_T_1018_mask) begin
      ram_header_src[ram_header_src_T_1018_addr] <= ram_header_src_T_1018_data;
    end
    if(ram_header_dst_T_1018_en & ram_header_dst_T_1018_mask) begin
      ram_header_dst[ram_header_dst_T_1018_addr] <= ram_header_dst_T_1018_data;
    end
    if(ram_payload_addr_beat_T_1018_en & ram_payload_addr_beat_T_1018_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1018_addr] <= ram_payload_addr_beat_T_1018_data;
    end
    if(ram_payload_addr_block_T_1018_en & ram_payload_addr_block_T_1018_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1018_addr] <= ram_payload_addr_block_T_1018_data;
    end
    if(ram_payload_client_xact_id_T_1018_en & ram_payload_client_xact_id_T_1018_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1018_addr] <= ram_payload_client_xact_id_T_1018_data;
    end
    if(ram_payload_voluntary_T_1018_en & ram_payload_voluntary_T_1018_mask) begin
      ram_payload_voluntary[ram_payload_voluntary_T_1018_addr] <= ram_payload_voluntary_T_1018_data;
    end
    if(ram_payload_r_type_T_1018_en & ram_payload_r_type_T_1018_mask) begin
      ram_payload_r_type[ram_payload_r_type_T_1018_addr] <= ram_payload_r_type_T_1018_data;
    end
    if(ram_payload_data_T_1018_en & ram_payload_data_T_1018_mask) begin
      ram_payload_data[ram_payload_data_T_1018_addr] <= ram_payload_data_T_1018_data;
    end
    if(reset) begin
      T_1010 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_1010 <= T_1133;
      end
    end
    if(reset) begin
      T_1012 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_1012 <= T_1138;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_3(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input   io_enq_bits_payload_client_xact_id,
  input  [1:0] io_enq_bits_payload_manager_xact_id,
  input   io_enq_bits_payload_is_builtin_type,
  input  [3:0] io_enq_bits_payload_g_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output  io_deq_bits_payload_client_xact_id,
  output [1:0] io_deq_bits_payload_manager_xact_id,
  output  io_deq_bits_payload_is_builtin_type,
  output [3:0] io_deq_bits_payload_g_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [1:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1144_data;
  wire  ram_header_src_T_1144_addr;
  wire  ram_header_src_T_1144_en;
  wire [1:0] ram_header_src_T_1018_data;
  wire  ram_header_src_T_1018_addr;
  wire  ram_header_src_T_1018_mask;
  wire  ram_header_src_T_1018_en;
  reg [1:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1144_data;
  wire  ram_header_dst_T_1144_addr;
  wire  ram_header_dst_T_1144_en;
  wire [1:0] ram_header_dst_T_1018_data;
  wire  ram_header_dst_T_1018_addr;
  wire  ram_header_dst_T_1018_mask;
  wire  ram_header_dst_T_1018_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1144_data;
  wire  ram_payload_addr_beat_T_1144_addr;
  wire  ram_payload_addr_beat_T_1144_en;
  wire [2:0] ram_payload_addr_beat_T_1018_data;
  wire  ram_payload_addr_beat_T_1018_addr;
  wire  ram_payload_addr_beat_T_1018_mask;
  wire  ram_payload_addr_beat_T_1018_en;
  reg  ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_3;
  wire  ram_payload_client_xact_id_T_1144_data;
  wire  ram_payload_client_xact_id_T_1144_addr;
  wire  ram_payload_client_xact_id_T_1144_en;
  wire  ram_payload_client_xact_id_T_1018_data;
  wire  ram_payload_client_xact_id_T_1018_addr;
  wire  ram_payload_client_xact_id_T_1018_mask;
  wire  ram_payload_client_xact_id_T_1018_en;
  reg [1:0] ram_payload_manager_xact_id [0:1];
  reg [31:0] GEN_4;
  wire [1:0] ram_payload_manager_xact_id_T_1144_data;
  wire  ram_payload_manager_xact_id_T_1144_addr;
  wire  ram_payload_manager_xact_id_T_1144_en;
  wire [1:0] ram_payload_manager_xact_id_T_1018_data;
  wire  ram_payload_manager_xact_id_T_1018_addr;
  wire  ram_payload_manager_xact_id_T_1018_mask;
  wire  ram_payload_manager_xact_id_T_1018_en;
  reg  ram_payload_is_builtin_type [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1144_data;
  wire  ram_payload_is_builtin_type_T_1144_addr;
  wire  ram_payload_is_builtin_type_T_1144_en;
  wire  ram_payload_is_builtin_type_T_1018_data;
  wire  ram_payload_is_builtin_type_T_1018_addr;
  wire  ram_payload_is_builtin_type_T_1018_mask;
  wire  ram_payload_is_builtin_type_T_1018_en;
  reg [3:0] ram_payload_g_type [0:1];
  reg [31:0] GEN_6;
  wire [3:0] ram_payload_g_type_T_1144_data;
  wire  ram_payload_g_type_T_1144_addr;
  wire  ram_payload_g_type_T_1144_en;
  wire [3:0] ram_payload_g_type_T_1018_data;
  wire  ram_payload_g_type_T_1018_addr;
  wire  ram_payload_g_type_T_1018_mask;
  wire  ram_payload_g_type_T_1018_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1144_data;
  wire  ram_payload_data_T_1144_addr;
  wire  ram_payload_data_T_1144_en;
  wire [63:0] ram_payload_data_T_1018_data;
  wire  ram_payload_data_T_1018_addr;
  wire  ram_payload_data_T_1018_mask;
  wire  ram_payload_data_T_1018_en;
  reg  T_1010;
  reg [31:0] GEN_8;
  reg  T_1012;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1015;
  wire  empty;
  wire  full;
  wire  T_1016;
  wire  do_enq;
  wire  T_1017;
  wire  do_deq;
  wire [1:0] T_1132;
  wire  T_1133;
  wire  GEN_19;
  wire [1:0] T_1137;
  wire  T_1138;
  wire  GEN_20;
  wire  T_1139;
  wire  GEN_21;
  wire  T_1141;
  wire  T_1143;
  wire [1:0] T_1255;
  wire  ptr_diff;
  wire  T_1256;
  wire [1:0] T_1257;
  assign io_enq_ready = T_1143;
  assign io_deq_valid = T_1141;
  assign io_deq_bits_header_src = ram_header_src_T_1144_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1144_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1144_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1144_data;
  assign io_deq_bits_payload_manager_xact_id = ram_payload_manager_xact_id_T_1144_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1144_data;
  assign io_deq_bits_payload_g_type = ram_payload_g_type_T_1144_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1144_data;
  assign io_count = T_1257;
  assign ram_header_src_T_1144_addr = T_1012;
  assign ram_header_src_T_1144_en = 1'h1;
  assign ram_header_src_T_1144_data = ram_header_src[ram_header_src_T_1144_addr];
  assign ram_header_src_T_1018_data = io_enq_bits_header_src;
  assign ram_header_src_T_1018_addr = T_1010;
  assign ram_header_src_T_1018_mask = do_enq;
  assign ram_header_src_T_1018_en = do_enq;
  assign ram_header_dst_T_1144_addr = T_1012;
  assign ram_header_dst_T_1144_en = 1'h1;
  assign ram_header_dst_T_1144_data = ram_header_dst[ram_header_dst_T_1144_addr];
  assign ram_header_dst_T_1018_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1018_addr = T_1010;
  assign ram_header_dst_T_1018_mask = do_enq;
  assign ram_header_dst_T_1018_en = do_enq;
  assign ram_payload_addr_beat_T_1144_addr = T_1012;
  assign ram_payload_addr_beat_T_1144_en = 1'h1;
  assign ram_payload_addr_beat_T_1144_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1144_addr];
  assign ram_payload_addr_beat_T_1018_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1018_addr = T_1010;
  assign ram_payload_addr_beat_T_1018_mask = do_enq;
  assign ram_payload_addr_beat_T_1018_en = do_enq;
  assign ram_payload_client_xact_id_T_1144_addr = T_1012;
  assign ram_payload_client_xact_id_T_1144_en = 1'h1;
  assign ram_payload_client_xact_id_T_1144_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1144_addr];
  assign ram_payload_client_xact_id_T_1018_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1018_addr = T_1010;
  assign ram_payload_client_xact_id_T_1018_mask = do_enq;
  assign ram_payload_client_xact_id_T_1018_en = do_enq;
  assign ram_payload_manager_xact_id_T_1144_addr = T_1012;
  assign ram_payload_manager_xact_id_T_1144_en = 1'h1;
  assign ram_payload_manager_xact_id_T_1144_data = ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1144_addr];
  assign ram_payload_manager_xact_id_T_1018_data = io_enq_bits_payload_manager_xact_id;
  assign ram_payload_manager_xact_id_T_1018_addr = T_1010;
  assign ram_payload_manager_xact_id_T_1018_mask = do_enq;
  assign ram_payload_manager_xact_id_T_1018_en = do_enq;
  assign ram_payload_is_builtin_type_T_1144_addr = T_1012;
  assign ram_payload_is_builtin_type_T_1144_en = 1'h1;
  assign ram_payload_is_builtin_type_T_1144_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1144_addr];
  assign ram_payload_is_builtin_type_T_1018_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1018_addr = T_1010;
  assign ram_payload_is_builtin_type_T_1018_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1018_en = do_enq;
  assign ram_payload_g_type_T_1144_addr = T_1012;
  assign ram_payload_g_type_T_1144_en = 1'h1;
  assign ram_payload_g_type_T_1144_data = ram_payload_g_type[ram_payload_g_type_T_1144_addr];
  assign ram_payload_g_type_T_1018_data = io_enq_bits_payload_g_type;
  assign ram_payload_g_type_T_1018_addr = T_1010;
  assign ram_payload_g_type_T_1018_mask = do_enq;
  assign ram_payload_g_type_T_1018_en = do_enq;
  assign ram_payload_data_T_1144_addr = T_1012;
  assign ram_payload_data_T_1144_en = 1'h1;
  assign ram_payload_data_T_1144_data = ram_payload_data[ram_payload_data_T_1144_addr];
  assign ram_payload_data_T_1018_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1018_addr = T_1010;
  assign ram_payload_data_T_1018_mask = do_enq;
  assign ram_payload_data_T_1018_en = do_enq;
  assign ptr_match = T_1010 == T_1012;
  assign T_1015 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1015;
  assign full = ptr_match & maybe_full;
  assign T_1016 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1016;
  assign T_1017 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1017;
  assign T_1132 = T_1010 + 1'h1;
  assign T_1133 = T_1132[0:0];
  assign GEN_19 = do_enq ? T_1133 : T_1010;
  assign T_1137 = T_1012 + 1'h1;
  assign T_1138 = T_1137[0:0];
  assign GEN_20 = do_deq ? T_1138 : T_1012;
  assign T_1139 = do_enq != do_deq;
  assign GEN_21 = T_1139 ? do_enq : maybe_full;
  assign T_1141 = empty == 1'h0;
  assign T_1143 = full == 1'h0;
  assign T_1255 = T_1010 - T_1012;
  assign ptr_diff = T_1255[0:0];
  assign T_1256 = maybe_full & ptr_match;
  assign T_1257 = {T_1256,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_manager_xact_id[initvar] = GEN_4[1:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_g_type[initvar] = GEN_6[3:0];
  `endif
  GEN_7 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  T_1010 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {1{$random}};
  T_1012 = GEN_9[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1018_en & ram_header_src_T_1018_mask) begin
      ram_header_src[ram_header_src_T_1018_addr] <= ram_header_src_T_1018_data;
    end
    if(ram_header_dst_T_1018_en & ram_header_dst_T_1018_mask) begin
      ram_header_dst[ram_header_dst_T_1018_addr] <= ram_header_dst_T_1018_data;
    end
    if(ram_payload_addr_beat_T_1018_en & ram_payload_addr_beat_T_1018_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1018_addr] <= ram_payload_addr_beat_T_1018_data;
    end
    if(ram_payload_client_xact_id_T_1018_en & ram_payload_client_xact_id_T_1018_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1018_addr] <= ram_payload_client_xact_id_T_1018_data;
    end
    if(ram_payload_manager_xact_id_T_1018_en & ram_payload_manager_xact_id_T_1018_mask) begin
      ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1018_addr] <= ram_payload_manager_xact_id_T_1018_data;
    end
    if(ram_payload_is_builtin_type_T_1018_en & ram_payload_is_builtin_type_T_1018_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1018_addr] <= ram_payload_is_builtin_type_T_1018_data;
    end
    if(ram_payload_g_type_T_1018_en & ram_payload_g_type_T_1018_mask) begin
      ram_payload_g_type[ram_payload_g_type_T_1018_addr] <= ram_payload_g_type_T_1018_data;
    end
    if(ram_payload_data_T_1018_en & ram_payload_data_T_1018_mask) begin
      ram_payload_data[ram_payload_data_T_1018_addr] <= ram_payload_data_T_1018_data;
    end
    if(reset) begin
      T_1010 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_1010 <= T_1133;
      end
    end
    if(reset) begin
      T_1012 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_1012 <= T_1138;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module TileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input   io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [10:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output  io_client_grant_bits_payload_client_xact_id,
  output [1:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [1:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input   io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output  io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [10:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input   io_manager_grant_bits_payload_client_xact_id,
  input  [1:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [1:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output  io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_4_clk;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [1:0] Queue_4_io_enq_bits_header_src;
  wire [1:0] Queue_4_io_enq_bits_header_dst;
  wire [25:0] Queue_4_io_enq_bits_payload_addr_block;
  wire  Queue_4_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_4_io_enq_bits_payload_addr_beat;
  wire  Queue_4_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_4_io_enq_bits_payload_a_type;
  wire [10:0] Queue_4_io_enq_bits_payload_union;
  wire [63:0] Queue_4_io_enq_bits_payload_data;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [1:0] Queue_4_io_deq_bits_header_src;
  wire [1:0] Queue_4_io_deq_bits_header_dst;
  wire [25:0] Queue_4_io_deq_bits_payload_addr_block;
  wire  Queue_4_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_4_io_deq_bits_payload_addr_beat;
  wire  Queue_4_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_4_io_deq_bits_payload_a_type;
  wire [10:0] Queue_4_io_deq_bits_payload_union;
  wire [63:0] Queue_4_io_deq_bits_payload_data;
  wire  Queue_4_io_count;
  wire  Queue_1_1_clk;
  wire  Queue_1_1_reset;
  wire  Queue_1_1_io_enq_ready;
  wire  Queue_1_1_io_enq_valid;
  wire [1:0] Queue_1_1_io_enq_bits_header_src;
  wire [1:0] Queue_1_1_io_enq_bits_header_dst;
  wire [25:0] Queue_1_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_1_1_io_enq_bits_payload_p_type;
  wire  Queue_1_1_io_deq_ready;
  wire  Queue_1_1_io_deq_valid;
  wire [1:0] Queue_1_1_io_deq_bits_header_src;
  wire [1:0] Queue_1_1_io_deq_bits_header_dst;
  wire [25:0] Queue_1_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_1_1_io_deq_bits_payload_p_type;
  wire  Queue_1_1_io_count;
  wire  Queue_2_1_clk;
  wire  Queue_2_1_reset;
  wire  Queue_2_1_io_enq_ready;
  wire  Queue_2_1_io_enq_valid;
  wire [1:0] Queue_2_1_io_enq_bits_header_src;
  wire [1:0] Queue_2_1_io_enq_bits_header_dst;
  wire [2:0] Queue_2_1_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_2_1_io_enq_bits_payload_addr_block;
  wire  Queue_2_1_io_enq_bits_payload_client_xact_id;
  wire  Queue_2_1_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_2_1_io_enq_bits_payload_r_type;
  wire [63:0] Queue_2_1_io_enq_bits_payload_data;
  wire  Queue_2_1_io_deq_ready;
  wire  Queue_2_1_io_deq_valid;
  wire [1:0] Queue_2_1_io_deq_bits_header_src;
  wire [1:0] Queue_2_1_io_deq_bits_header_dst;
  wire [2:0] Queue_2_1_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_2_1_io_deq_bits_payload_addr_block;
  wire  Queue_2_1_io_deq_bits_payload_client_xact_id;
  wire  Queue_2_1_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_2_1_io_deq_bits_payload_r_type;
  wire [63:0] Queue_2_1_io_deq_bits_payload_data;
  wire [1:0] Queue_2_1_io_count;
  wire  Queue_3_1_clk;
  wire  Queue_3_1_reset;
  wire  Queue_3_1_io_enq_ready;
  wire  Queue_3_1_io_enq_valid;
  wire [1:0] Queue_3_1_io_enq_bits_header_src;
  wire [1:0] Queue_3_1_io_enq_bits_header_dst;
  wire [2:0] Queue_3_1_io_enq_bits_payload_addr_beat;
  wire  Queue_3_1_io_enq_bits_payload_client_xact_id;
  wire [1:0] Queue_3_1_io_enq_bits_payload_manager_xact_id;
  wire  Queue_3_1_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_3_1_io_enq_bits_payload_g_type;
  wire [63:0] Queue_3_1_io_enq_bits_payload_data;
  wire  Queue_3_1_io_deq_ready;
  wire  Queue_3_1_io_deq_valid;
  wire [1:0] Queue_3_1_io_deq_bits_header_src;
  wire [1:0] Queue_3_1_io_deq_bits_header_dst;
  wire [2:0] Queue_3_1_io_deq_bits_payload_addr_beat;
  wire  Queue_3_1_io_deq_bits_payload_client_xact_id;
  wire [1:0] Queue_3_1_io_deq_bits_payload_manager_xact_id;
  wire  Queue_3_1_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_3_1_io_deq_bits_payload_g_type;
  wire [63:0] Queue_3_1_io_deq_bits_payload_data;
  wire [1:0] Queue_3_1_io_count;
  Queue Queue_4 (
    .clk(Queue_4_clk),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_header_src(Queue_4_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_4_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_4_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_4_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_4_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_4_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_4_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_4_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_4_io_enq_bits_payload_data),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_header_src(Queue_4_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_4_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_4_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_4_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_4_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_4_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_4_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_4_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_4_io_deq_bits_payload_data),
    .io_count(Queue_4_io_count)
  );
  Queue_1 Queue_1_1 (
    .clk(Queue_1_1_clk),
    .reset(Queue_1_1_reset),
    .io_enq_ready(Queue_1_1_io_enq_ready),
    .io_enq_valid(Queue_1_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_1_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_1_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_1_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_1_1_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_1_1_io_deq_ready),
    .io_deq_valid(Queue_1_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_1_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_1_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_1_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_1_1_io_deq_bits_payload_p_type),
    .io_count(Queue_1_1_io_count)
  );
  Queue_2 Queue_2_1 (
    .clk(Queue_2_1_clk),
    .reset(Queue_2_1_reset),
    .io_enq_ready(Queue_2_1_io_enq_ready),
    .io_enq_valid(Queue_2_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_2_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_2_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_2_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_2_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_2_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_2_1_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_2_1_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_2_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_2_1_io_deq_ready),
    .io_deq_valid(Queue_2_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_2_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_2_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_2_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_2_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_2_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_2_1_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_2_1_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_2_1_io_deq_bits_payload_data),
    .io_count(Queue_2_1_io_count)
  );
  Queue_3 Queue_3_1 (
    .clk(Queue_3_1_clk),
    .reset(Queue_3_1_reset),
    .io_enq_ready(Queue_3_1_io_enq_ready),
    .io_enq_valid(Queue_3_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_3_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_3_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_3_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_3_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_3_1_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_3_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_3_1_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_3_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_3_1_io_deq_ready),
    .io_deq_valid(Queue_3_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_3_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_3_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_3_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_3_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_3_1_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_3_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_3_1_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_3_1_io_deq_bits_payload_data),
    .io_count(Queue_3_1_io_count)
  );
  assign io_client_acquire_ready = Queue_4_io_enq_ready;
  assign io_client_grant_valid = Queue_3_1_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_3_1_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_3_1_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_3_1_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_3_1_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_3_1_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_3_1_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_3_1_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_3_1_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_1_1_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_1_1_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_1_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_1_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_1_1_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_2_1_io_enq_ready;
  assign io_manager_acquire_valid = Queue_4_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_4_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_4_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_4_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_4_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_4_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_4_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_4_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_4_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_4_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_3_1_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_1_1_io_enq_ready;
  assign io_manager_release_valid = Queue_2_1_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_2_1_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_2_1_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_2_1_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_2_1_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_2_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_2_1_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_2_1_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_2_1_io_deq_bits_payload_data;
  assign Queue_4_clk = clk;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = io_client_acquire_valid;
  assign Queue_4_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_4_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_4_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_4_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_4_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_4_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_4_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_4_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_4_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_4_io_deq_ready = io_manager_acquire_ready;
  assign Queue_1_1_clk = clk;
  assign Queue_1_1_reset = reset;
  assign Queue_1_1_io_enq_valid = io_manager_probe_valid;
  assign Queue_1_1_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_1_1_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_1_1_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_1_1_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_1_1_io_deq_ready = io_client_probe_ready;
  assign Queue_2_1_clk = clk;
  assign Queue_2_1_reset = reset;
  assign Queue_2_1_io_enq_valid = io_client_release_valid;
  assign Queue_2_1_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_2_1_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_2_1_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_2_1_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_2_1_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_2_1_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_2_1_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_2_1_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_2_1_io_deq_ready = io_manager_release_ready;
  assign Queue_3_1_clk = clk;
  assign Queue_3_1_reset = reset;
  assign Queue_3_1_io_enq_valid = io_manager_grant_valid;
  assign Queue_3_1_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_3_1_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_3_1_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_3_1_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_3_1_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_3_1_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_3_1_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_3_1_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_3_1_io_deq_ready = io_client_grant_ready;
endmodule
module ClientTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input   io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [10:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [25:0] io_client_probe_bits_addr_block,
  output [1:0] io_client_probe_bits_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [2:0] io_client_release_bits_addr_beat,
  input  [25:0] io_client_release_bits_addr_block,
  input   io_client_release_bits_client_xact_id,
  input   io_client_release_bits_voluntary,
  input  [2:0] io_client_release_bits_r_type,
  input  [63:0] io_client_release_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output  io_client_grant_bits_client_xact_id,
  output [1:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  output  io_client_grant_bits_manager_id,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_manager_xact_id,
  input   io_client_finish_bits_manager_id,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [1:0] io_network_acquire_bits_header_src,
  output [1:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output  io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [10:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [1:0] io_network_grant_bits_header_src,
  input  [1:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input   io_network_grant_bits_payload_client_xact_id,
  input  [1:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [1:0] io_network_finish_bits_header_src,
  output [1:0] io_network_finish_bits_header_dst,
  output [1:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [1:0] io_network_probe_bits_header_src,
  input  [1:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [1:0] io_network_release_bits_header_src,
  output [1:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output  io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [1:0] acq_with_header_bits_header_src;
  wire [1:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire  acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [10:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_3894;
  wire  T_3896;
  wire  T_3898;
  wire  T_3899;
  wire  T_3902;
  wire  rel_with_header_ready;
  wire  rel_with_header_valid;
  wire [1:0] rel_with_header_bits_header_src;
  wire [1:0] rel_with_header_bits_header_dst;
  wire [2:0] rel_with_header_bits_payload_addr_beat;
  wire [25:0] rel_with_header_bits_payload_addr_block;
  wire  rel_with_header_bits_payload_client_xact_id;
  wire  rel_with_header_bits_payload_voluntary;
  wire [2:0] rel_with_header_bits_payload_r_type;
  wire [63:0] rel_with_header_bits_payload_data;
  wire [31:0] GEN_1;
  wire [31:0] T_4464;
  wire  T_4466;
  wire  T_4468;
  wire  T_4469;
  wire  T_4472;
  wire  fin_with_header_ready;
  wire  fin_with_header_valid;
  wire [1:0] fin_with_header_bits_header_src;
  wire [1:0] fin_with_header_bits_header_dst;
  wire [1:0] fin_with_header_bits_payload_manager_xact_id;
  wire  fin_with_header_bits_payload_manager_id;
  wire  prb_without_header_ready;
  wire  prb_without_header_valid;
  wire [25:0] prb_without_header_bits_addr_block;
  wire [1:0] prb_without_header_bits_p_type;
  wire  gnt_without_header_ready;
  wire  gnt_without_header_valid;
  wire [2:0] gnt_without_header_bits_addr_beat;
  wire  gnt_without_header_bits_client_xact_id;
  wire [1:0] gnt_without_header_bits_manager_xact_id;
  wire  gnt_without_header_bits_is_builtin_type;
  wire [3:0] gnt_without_header_bits_g_type;
  wire [63:0] gnt_without_header_bits_data;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_probe_valid = prb_without_header_valid;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign io_client_release_ready = rel_with_header_ready;
  assign io_client_grant_valid = gnt_without_header_valid;
  assign io_client_grant_bits_addr_beat = gnt_without_header_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = gnt_without_header_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = gnt_without_header_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = gnt_without_header_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = gnt_without_header_bits_g_type;
  assign io_client_grant_bits_data = gnt_without_header_bits_data;
  assign io_client_grant_bits_manager_id = io_network_grant_bits_header_src[0];
  assign io_client_finish_ready = fin_with_header_ready;
  assign io_network_acquire_valid = acq_with_header_valid;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = gnt_without_header_ready;
  assign io_network_finish_valid = fin_with_header_valid;
  assign io_network_finish_bits_header_src = fin_with_header_bits_header_src;
  assign io_network_finish_bits_header_dst = fin_with_header_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = fin_with_header_bits_payload_manager_xact_id;
  assign io_network_probe_ready = prb_without_header_ready;
  assign io_network_release_valid = rel_with_header_valid;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign acq_with_header_ready = io_network_acquire_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = 2'h0;
  assign acq_with_header_bits_header_dst = {{1'd0}, T_3902};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_3894 = GEN_0 << 6;
  assign T_3896 = 32'h80000000 <= T_3894;
  assign T_3898 = T_3894 < 32'h90000000;
  assign T_3899 = T_3896 & T_3898;
  assign T_3902 = T_3899 ? 1'h0 : 1'h1;
  assign rel_with_header_ready = io_network_release_ready;
  assign rel_with_header_valid = io_client_release_valid;
  assign rel_with_header_bits_header_src = 2'h0;
  assign rel_with_header_bits_header_dst = {{1'd0}, T_4472};
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign GEN_1 = {{6'd0}, io_client_release_bits_addr_block};
  assign T_4464 = GEN_1 << 6;
  assign T_4466 = 32'h80000000 <= T_4464;
  assign T_4468 = T_4464 < 32'h90000000;
  assign T_4469 = T_4466 & T_4468;
  assign T_4472 = T_4469 ? 1'h0 : 1'h1;
  assign fin_with_header_ready = io_network_finish_ready;
  assign fin_with_header_valid = io_client_finish_valid;
  assign fin_with_header_bits_header_src = 2'h0;
  assign fin_with_header_bits_header_dst = {{1'd0}, io_client_finish_bits_manager_id};
  assign fin_with_header_bits_payload_manager_xact_id = io_client_finish_bits_manager_xact_id;
  assign fin_with_header_bits_payload_manager_id = io_client_finish_bits_manager_id;
  assign prb_without_header_ready = io_client_probe_ready;
  assign prb_without_header_valid = io_network_probe_valid;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign gnt_without_header_ready = io_client_grant_ready;
  assign gnt_without_header_valid = io_network_grant_valid;
  assign gnt_without_header_bits_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign gnt_without_header_bits_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign gnt_without_header_bits_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign gnt_without_header_bits_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign gnt_without_header_bits_g_type = io_network_grant_bits_payload_g_type;
  assign gnt_without_header_bits_data = io_network_grant_bits_payload_data;
endmodule
module TileLinkEnqueuer_1(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input   io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [10:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output  io_client_grant_bits_payload_client_xact_id,
  output [1:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [1:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input   io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output  io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [10:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input   io_manager_grant_bits_payload_client_xact_id,
  input  [1:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [1:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output  io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_4_1_clk;
  wire  Queue_4_1_reset;
  wire  Queue_4_1_io_enq_ready;
  wire  Queue_4_1_io_enq_valid;
  wire [1:0] Queue_4_1_io_enq_bits_header_src;
  wire [1:0] Queue_4_1_io_enq_bits_header_dst;
  wire [25:0] Queue_4_1_io_enq_bits_payload_addr_block;
  wire  Queue_4_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_4_1_io_enq_bits_payload_addr_beat;
  wire  Queue_4_1_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_4_1_io_enq_bits_payload_a_type;
  wire [10:0] Queue_4_1_io_enq_bits_payload_union;
  wire [63:0] Queue_4_1_io_enq_bits_payload_data;
  wire  Queue_4_1_io_deq_ready;
  wire  Queue_4_1_io_deq_valid;
  wire [1:0] Queue_4_1_io_deq_bits_header_src;
  wire [1:0] Queue_4_1_io_deq_bits_header_dst;
  wire [25:0] Queue_4_1_io_deq_bits_payload_addr_block;
  wire  Queue_4_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_4_1_io_deq_bits_payload_addr_beat;
  wire  Queue_4_1_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_4_1_io_deq_bits_payload_a_type;
  wire [10:0] Queue_4_1_io_deq_bits_payload_union;
  wire [63:0] Queue_4_1_io_deq_bits_payload_data;
  wire  Queue_4_1_io_count;
  wire  Queue_5_1_clk;
  wire  Queue_5_1_reset;
  wire  Queue_5_1_io_enq_ready;
  wire  Queue_5_1_io_enq_valid;
  wire [1:0] Queue_5_1_io_enq_bits_header_src;
  wire [1:0] Queue_5_1_io_enq_bits_header_dst;
  wire [25:0] Queue_5_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_5_1_io_enq_bits_payload_p_type;
  wire  Queue_5_1_io_deq_ready;
  wire  Queue_5_1_io_deq_valid;
  wire [1:0] Queue_5_1_io_deq_bits_header_src;
  wire [1:0] Queue_5_1_io_deq_bits_header_dst;
  wire [25:0] Queue_5_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_5_1_io_deq_bits_payload_p_type;
  wire  Queue_5_1_io_count;
  wire  Queue_6_1_clk;
  wire  Queue_6_1_reset;
  wire  Queue_6_1_io_enq_ready;
  wire  Queue_6_1_io_enq_valid;
  wire [1:0] Queue_6_1_io_enq_bits_header_src;
  wire [1:0] Queue_6_1_io_enq_bits_header_dst;
  wire [2:0] Queue_6_1_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_6_1_io_enq_bits_payload_addr_block;
  wire  Queue_6_1_io_enq_bits_payload_client_xact_id;
  wire  Queue_6_1_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_6_1_io_enq_bits_payload_r_type;
  wire [63:0] Queue_6_1_io_enq_bits_payload_data;
  wire  Queue_6_1_io_deq_ready;
  wire  Queue_6_1_io_deq_valid;
  wire [1:0] Queue_6_1_io_deq_bits_header_src;
  wire [1:0] Queue_6_1_io_deq_bits_header_dst;
  wire [2:0] Queue_6_1_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_6_1_io_deq_bits_payload_addr_block;
  wire  Queue_6_1_io_deq_bits_payload_client_xact_id;
  wire  Queue_6_1_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_6_1_io_deq_bits_payload_r_type;
  wire [63:0] Queue_6_1_io_deq_bits_payload_data;
  wire [1:0] Queue_6_1_io_count;
  wire  Queue_7_1_clk;
  wire  Queue_7_1_reset;
  wire  Queue_7_1_io_enq_ready;
  wire  Queue_7_1_io_enq_valid;
  wire [1:0] Queue_7_1_io_enq_bits_header_src;
  wire [1:0] Queue_7_1_io_enq_bits_header_dst;
  wire [2:0] Queue_7_1_io_enq_bits_payload_addr_beat;
  wire  Queue_7_1_io_enq_bits_payload_client_xact_id;
  wire [1:0] Queue_7_1_io_enq_bits_payload_manager_xact_id;
  wire  Queue_7_1_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_7_1_io_enq_bits_payload_g_type;
  wire [63:0] Queue_7_1_io_enq_bits_payload_data;
  wire  Queue_7_1_io_deq_ready;
  wire  Queue_7_1_io_deq_valid;
  wire [1:0] Queue_7_1_io_deq_bits_header_src;
  wire [1:0] Queue_7_1_io_deq_bits_header_dst;
  wire [2:0] Queue_7_1_io_deq_bits_payload_addr_beat;
  wire  Queue_7_1_io_deq_bits_payload_client_xact_id;
  wire [1:0] Queue_7_1_io_deq_bits_payload_manager_xact_id;
  wire  Queue_7_1_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_7_1_io_deq_bits_payload_g_type;
  wire [63:0] Queue_7_1_io_deq_bits_payload_data;
  wire [1:0] Queue_7_1_io_count;
  Queue Queue_4_1 (
    .clk(Queue_4_1_clk),
    .reset(Queue_4_1_reset),
    .io_enq_ready(Queue_4_1_io_enq_ready),
    .io_enq_valid(Queue_4_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_4_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_4_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_4_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_4_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_4_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_4_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_4_1_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_4_1_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_4_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_4_1_io_deq_ready),
    .io_deq_valid(Queue_4_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_4_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_4_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_4_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_4_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_4_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_4_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_4_1_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_4_1_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_4_1_io_deq_bits_payload_data),
    .io_count(Queue_4_1_io_count)
  );
  Queue_1 Queue_5_1 (
    .clk(Queue_5_1_clk),
    .reset(Queue_5_1_reset),
    .io_enq_ready(Queue_5_1_io_enq_ready),
    .io_enq_valid(Queue_5_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_5_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_5_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_5_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_5_1_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_5_1_io_deq_ready),
    .io_deq_valid(Queue_5_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_5_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_5_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_5_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_5_1_io_deq_bits_payload_p_type),
    .io_count(Queue_5_1_io_count)
  );
  Queue_2 Queue_6_1 (
    .clk(Queue_6_1_clk),
    .reset(Queue_6_1_reset),
    .io_enq_ready(Queue_6_1_io_enq_ready),
    .io_enq_valid(Queue_6_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_6_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_6_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_6_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_6_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_6_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_6_1_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_6_1_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_6_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_6_1_io_deq_ready),
    .io_deq_valid(Queue_6_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_6_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_6_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_6_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_6_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_6_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_6_1_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_6_1_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_6_1_io_deq_bits_payload_data),
    .io_count(Queue_6_1_io_count)
  );
  Queue_3 Queue_7_1 (
    .clk(Queue_7_1_clk),
    .reset(Queue_7_1_reset),
    .io_enq_ready(Queue_7_1_io_enq_ready),
    .io_enq_valid(Queue_7_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_7_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_7_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_7_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_7_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_7_1_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_7_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_7_1_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_7_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_7_1_io_deq_ready),
    .io_deq_valid(Queue_7_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_7_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_7_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_7_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_7_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_7_1_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_7_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_7_1_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_7_1_io_deq_bits_payload_data),
    .io_count(Queue_7_1_io_count)
  );
  assign io_client_acquire_ready = Queue_4_1_io_enq_ready;
  assign io_client_grant_valid = Queue_7_1_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_7_1_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_7_1_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_7_1_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_7_1_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_7_1_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_7_1_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_7_1_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_7_1_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_5_1_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_5_1_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_5_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_5_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_5_1_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_6_1_io_enq_ready;
  assign io_manager_acquire_valid = Queue_4_1_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_4_1_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_4_1_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_4_1_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_4_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_4_1_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_4_1_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_4_1_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_4_1_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_4_1_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_7_1_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_5_1_io_enq_ready;
  assign io_manager_release_valid = Queue_6_1_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_6_1_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_6_1_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_6_1_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_6_1_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_6_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_6_1_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_6_1_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_6_1_io_deq_bits_payload_data;
  assign Queue_4_1_clk = clk;
  assign Queue_4_1_reset = reset;
  assign Queue_4_1_io_enq_valid = io_client_acquire_valid;
  assign Queue_4_1_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_4_1_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_4_1_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_4_1_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_4_1_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_4_1_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_4_1_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_4_1_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_4_1_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_4_1_io_deq_ready = io_manager_acquire_ready;
  assign Queue_5_1_clk = clk;
  assign Queue_5_1_reset = reset;
  assign Queue_5_1_io_enq_valid = io_manager_probe_valid;
  assign Queue_5_1_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_5_1_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_5_1_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_5_1_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_5_1_io_deq_ready = io_client_probe_ready;
  assign Queue_6_1_clk = clk;
  assign Queue_6_1_reset = reset;
  assign Queue_6_1_io_enq_valid = io_client_release_valid;
  assign Queue_6_1_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_6_1_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_6_1_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_6_1_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_6_1_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_6_1_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_6_1_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_6_1_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_6_1_io_deq_ready = io_manager_release_ready;
  assign Queue_7_1_clk = clk;
  assign Queue_7_1_reset = reset;
  assign Queue_7_1_io_enq_valid = io_manager_grant_valid;
  assign Queue_7_1_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_7_1_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_7_1_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_7_1_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_7_1_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_7_1_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_7_1_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_7_1_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_7_1_io_deq_ready = io_client_grant_ready;
endmodule
module FinishQueue_1(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output [1:0] io_count
);
  reg [1:0] ram_manager_xact_id [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_manager_xact_id_T_264_data;
  wire  ram_manager_xact_id_T_264_addr;
  wire  ram_manager_xact_id_T_264_en;
  wire [1:0] ram_manager_xact_id_T_226_data;
  wire  ram_manager_xact_id_T_226_addr;
  wire  ram_manager_xact_id_T_226_mask;
  wire  ram_manager_xact_id_T_226_en;
  reg  ram_manager_id [0:1];
  reg [31:0] GEN_1;
  wire  ram_manager_id_T_264_data;
  wire  ram_manager_id_T_264_addr;
  wire  ram_manager_id_T_264_en;
  wire  ram_manager_id_T_226_data;
  wire  ram_manager_id_T_226_addr;
  wire  ram_manager_id_T_226_mask;
  wire  ram_manager_id_T_226_en;
  reg  T_218;
  reg [31:0] GEN_2;
  reg  T_220;
  reg [31:0] GEN_3;
  reg  maybe_full;
  reg [31:0] GEN_4;
  wire  ptr_match;
  wire  T_223;
  wire  empty;
  wire  full;
  wire  T_224;
  wire  do_enq;
  wire  T_225;
  wire  do_deq;
  wire [1:0] T_252;
  wire  T_253;
  wire  GEN_7;
  wire [1:0] T_257;
  wire  T_258;
  wire  GEN_8;
  wire  T_259;
  wire  GEN_9;
  wire  T_261;
  wire  T_263;
  wire [1:0] T_287;
  wire  ptr_diff;
  wire  T_288;
  wire [1:0] T_289;
  assign io_enq_ready = T_263;
  assign io_deq_valid = T_261;
  assign io_deq_bits_manager_xact_id = ram_manager_xact_id_T_264_data;
  assign io_deq_bits_manager_id = ram_manager_id_T_264_data;
  assign io_count = T_289;
  assign ram_manager_xact_id_T_264_addr = T_220;
  assign ram_manager_xact_id_T_264_en = 1'h1;
  assign ram_manager_xact_id_T_264_data = ram_manager_xact_id[ram_manager_xact_id_T_264_addr];
  assign ram_manager_xact_id_T_226_data = io_enq_bits_manager_xact_id;
  assign ram_manager_xact_id_T_226_addr = T_218;
  assign ram_manager_xact_id_T_226_mask = do_enq;
  assign ram_manager_xact_id_T_226_en = do_enq;
  assign ram_manager_id_T_264_addr = T_220;
  assign ram_manager_id_T_264_en = 1'h1;
  assign ram_manager_id_T_264_data = ram_manager_id[ram_manager_id_T_264_addr];
  assign ram_manager_id_T_226_data = io_enq_bits_manager_id;
  assign ram_manager_id_T_226_addr = T_218;
  assign ram_manager_id_T_226_mask = do_enq;
  assign ram_manager_id_T_226_en = do_enq;
  assign ptr_match = T_218 == T_220;
  assign T_223 = maybe_full == 1'h0;
  assign empty = ptr_match & T_223;
  assign full = ptr_match & maybe_full;
  assign T_224 = io_enq_ready & io_enq_valid;
  assign do_enq = T_224;
  assign T_225 = io_deq_ready & io_deq_valid;
  assign do_deq = T_225;
  assign T_252 = T_218 + 1'h1;
  assign T_253 = T_252[0:0];
  assign GEN_7 = do_enq ? T_253 : T_218;
  assign T_257 = T_220 + 1'h1;
  assign T_258 = T_257[0:0];
  assign GEN_8 = do_deq ? T_258 : T_220;
  assign T_259 = do_enq != do_deq;
  assign GEN_9 = T_259 ? do_enq : maybe_full;
  assign T_261 = empty == 1'h0;
  assign T_263 = full == 1'h0;
  assign T_287 = T_218 - T_220;
  assign ptr_diff = T_287[0:0];
  assign T_288 = maybe_full & ptr_match;
  assign T_289 = {T_288,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_manager_xact_id[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_manager_id[initvar] = GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_218 = GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  T_220 = GEN_3[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {1{$random}};
  maybe_full = GEN_4[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_manager_xact_id_T_226_en & ram_manager_xact_id_T_226_mask) begin
      ram_manager_xact_id[ram_manager_xact_id_T_226_addr] <= ram_manager_xact_id_T_226_data;
    end
    if(ram_manager_id_T_226_en & ram_manager_id_T_226_mask) begin
      ram_manager_id[ram_manager_id_T_226_addr] <= ram_manager_id_T_226_data;
    end
    if(reset) begin
      T_218 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_218 <= T_253;
      end
    end
    if(reset) begin
      T_220 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_220 <= T_258;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_259) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module FinishUnit(
  input   clk,
  input   reset,
  output  io_grant_ready,
  input   io_grant_valid,
  input  [1:0] io_grant_bits_header_src,
  input  [1:0] io_grant_bits_header_dst,
  input  [2:0] io_grant_bits_payload_addr_beat,
  input   io_grant_bits_payload_client_xact_id,
  input  [1:0] io_grant_bits_payload_manager_xact_id,
  input   io_grant_bits_payload_is_builtin_type,
  input  [3:0] io_grant_bits_payload_g_type,
  input  [63:0] io_grant_bits_payload_data,
  input   io_refill_ready,
  output  io_refill_valid,
  output [2:0] io_refill_bits_addr_beat,
  output  io_refill_bits_client_xact_id,
  output [1:0] io_refill_bits_manager_xact_id,
  output  io_refill_bits_is_builtin_type,
  output [3:0] io_refill_bits_g_type,
  output [63:0] io_refill_bits_data,
  input   io_finish_ready,
  output  io_finish_valid,
  output [1:0] io_finish_bits_header_src,
  output [1:0] io_finish_bits_header_dst,
  output [1:0] io_finish_bits_payload_manager_xact_id,
  output  io_ready
);
  wire  T_1035;
  wire [2:0] T_1044_0;
  wire [3:0] GEN_1;
  wire  T_1046;
  wire  T_1047;
  wire  T_1048;
  wire  T_1050;
  reg [2:0] T_1052;
  reg [31:0] GEN_3;
  wire  T_1054;
  wire [3:0] T_1056;
  wire [2:0] T_1057;
  wire [2:0] GEN_0;
  wire  T_1058;
  wire  T_1060;
  wire  FinishQueue_1_1_clk;
  wire  FinishQueue_1_1_reset;
  wire  FinishQueue_1_1_io_enq_ready;
  wire  FinishQueue_1_1_io_enq_valid;
  wire [1:0] FinishQueue_1_1_io_enq_bits_manager_xact_id;
  wire  FinishQueue_1_1_io_enq_bits_manager_id;
  wire  FinishQueue_1_1_io_deq_ready;
  wire  FinishQueue_1_1_io_deq_valid;
  wire [1:0] FinishQueue_1_1_io_deq_bits_manager_xact_id;
  wire  FinishQueue_1_1_io_deq_bits_manager_id;
  wire [1:0] FinishQueue_1_1_io_count;
  wire  T_1090;
  wire  T_1092;
  wire  T_1094;
  wire [2:0] T_1102_0;
  wire [3:0] GEN_2;
  wire  T_1104;
  wire  T_1106;
  wire  T_1109;
  wire  T_1110;
  wire  T_1111;
  wire [1:0] T_1134_manager_xact_id;
  wire  T_1167;
  wire  T_1168;
  wire  T_1169;
  wire  T_1182;
  FinishQueue_1 FinishQueue_1_1 (
    .clk(FinishQueue_1_1_clk),
    .reset(FinishQueue_1_1_reset),
    .io_enq_ready(FinishQueue_1_1_io_enq_ready),
    .io_enq_valid(FinishQueue_1_1_io_enq_valid),
    .io_enq_bits_manager_xact_id(FinishQueue_1_1_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(FinishQueue_1_1_io_enq_bits_manager_id),
    .io_deq_ready(FinishQueue_1_1_io_deq_ready),
    .io_deq_valid(FinishQueue_1_1_io_deq_valid),
    .io_deq_bits_manager_xact_id(FinishQueue_1_1_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(FinishQueue_1_1_io_deq_bits_manager_id),
    .io_count(FinishQueue_1_1_io_count)
  );
  assign io_grant_ready = T_1182;
  assign io_refill_valid = T_1169;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_finish_valid = FinishQueue_1_1_io_deq_valid;
  assign io_finish_bits_header_src = 2'h1;
  assign io_finish_bits_header_dst = {{1'd0}, FinishQueue_1_1_io_deq_bits_manager_id};
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_1_1_io_deq_bits_manager_xact_id;
  assign io_ready = FinishQueue_1_1_io_enq_ready;
  assign T_1035 = io_grant_ready & io_grant_valid;
  assign T_1044_0 = 3'h5;
  assign GEN_1 = {{1'd0}, T_1044_0};
  assign T_1046 = io_grant_bits_payload_g_type == GEN_1;
  assign T_1047 = io_grant_bits_payload_g_type == 4'h0;
  assign T_1048 = io_grant_bits_payload_is_builtin_type ? T_1046 : T_1047;
  assign T_1050 = T_1035 & T_1048;
  assign T_1054 = T_1052 == 3'h7;
  assign T_1056 = T_1052 + 3'h1;
  assign T_1057 = T_1056[2:0];
  assign GEN_0 = T_1050 ? T_1057 : T_1052;
  assign T_1058 = T_1050 & T_1054;
  assign T_1060 = T_1048 ? T_1058 : T_1035;
  assign FinishQueue_1_1_clk = clk;
  assign FinishQueue_1_1_reset = reset;
  assign FinishQueue_1_1_io_enq_valid = T_1111;
  assign FinishQueue_1_1_io_enq_bits_manager_xact_id = T_1134_manager_xact_id;
  assign FinishQueue_1_1_io_enq_bits_manager_id = io_grant_bits_header_src[0];
  assign FinishQueue_1_1_io_deq_ready = io_finish_ready;
  assign T_1090 = io_grant_bits_payload_is_builtin_type & T_1047;
  assign T_1092 = T_1090 == 1'h0;
  assign T_1094 = T_1035 & T_1092;
  assign T_1102_0 = 3'h5;
  assign GEN_2 = {{1'd0}, T_1102_0};
  assign T_1104 = io_grant_bits_payload_g_type == GEN_2;
  assign T_1106 = io_grant_bits_payload_is_builtin_type ? T_1104 : T_1047;
  assign T_1109 = T_1106 == 1'h0;
  assign T_1110 = T_1109 | T_1060;
  assign T_1111 = T_1094 & T_1110;
  assign T_1134_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign T_1167 = T_1092 == 1'h0;
  assign T_1168 = FinishQueue_1_1_io_enq_ready | T_1167;
  assign T_1169 = T_1168 & io_grant_valid;
  assign T_1182 = T_1168 & io_refill_ready;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  T_1052 = GEN_3[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1052 <= 3'h0;
    end else begin
      if(T_1050) begin
        T_1052 <= T_1057;
      end
    end
  end
endmodule
module ClientUncachedTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input   io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [10:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output  io_client_grant_bits_client_xact_id,
  output [1:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [1:0] io_network_acquire_bits_header_src,
  output [1:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output  io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [10:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [1:0] io_network_grant_bits_header_src,
  input  [1:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input   io_network_grant_bits_payload_client_xact_id,
  input  [1:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [1:0] io_network_finish_bits_header_src,
  output [1:0] io_network_finish_bits_header_dst,
  output [1:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [1:0] io_network_probe_bits_header_src,
  input  [1:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [1:0] io_network_release_bits_header_src,
  output [1:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output  io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  finisher_clk;
  wire  finisher_reset;
  wire  finisher_io_grant_ready;
  wire  finisher_io_grant_valid;
  wire [1:0] finisher_io_grant_bits_header_src;
  wire [1:0] finisher_io_grant_bits_header_dst;
  wire [2:0] finisher_io_grant_bits_payload_addr_beat;
  wire  finisher_io_grant_bits_payload_client_xact_id;
  wire [1:0] finisher_io_grant_bits_payload_manager_xact_id;
  wire  finisher_io_grant_bits_payload_is_builtin_type;
  wire [3:0] finisher_io_grant_bits_payload_g_type;
  wire [63:0] finisher_io_grant_bits_payload_data;
  wire  finisher_io_refill_ready;
  wire  finisher_io_refill_valid;
  wire [2:0] finisher_io_refill_bits_addr_beat;
  wire  finisher_io_refill_bits_client_xact_id;
  wire [1:0] finisher_io_refill_bits_manager_xact_id;
  wire  finisher_io_refill_bits_is_builtin_type;
  wire [3:0] finisher_io_refill_bits_g_type;
  wire [63:0] finisher_io_refill_bits_data;
  wire  finisher_io_finish_ready;
  wire  finisher_io_finish_valid;
  wire [1:0] finisher_io_finish_bits_header_src;
  wire [1:0] finisher_io_finish_bits_header_dst;
  wire [1:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire  finisher_io_ready;
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [1:0] acq_with_header_bits_header_src;
  wire [1:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire  acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [10:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_3330;
  wire  T_3332;
  wire  T_3334;
  wire  T_3335;
  wire  T_3338;
  wire  T_3339;
  wire  T_3340;
  wire [1:0] GEN_1;
  reg [31:0] GEN_9;
  wire [1:0] GEN_2;
  reg [31:0] GEN_10;
  wire [2:0] GEN_3;
  reg [31:0] GEN_11;
  wire [25:0] GEN_4;
  reg [31:0] GEN_12;
  wire  GEN_5;
  reg [31:0] GEN_13;
  wire  GEN_6;
  reg [31:0] GEN_14;
  wire [2:0] GEN_7;
  reg [31:0] GEN_15;
  wire [63:0] GEN_8;
  reg [63:0] GEN_16;
  FinishUnit finisher (
    .clk(finisher_clk),
    .reset(finisher_reset),
    .io_grant_ready(finisher_io_grant_ready),
    .io_grant_valid(finisher_io_grant_valid),
    .io_grant_bits_header_src(finisher_io_grant_bits_header_src),
    .io_grant_bits_header_dst(finisher_io_grant_bits_header_dst),
    .io_grant_bits_payload_addr_beat(finisher_io_grant_bits_payload_addr_beat),
    .io_grant_bits_payload_client_xact_id(finisher_io_grant_bits_payload_client_xact_id),
    .io_grant_bits_payload_manager_xact_id(finisher_io_grant_bits_payload_manager_xact_id),
    .io_grant_bits_payload_is_builtin_type(finisher_io_grant_bits_payload_is_builtin_type),
    .io_grant_bits_payload_g_type(finisher_io_grant_bits_payload_g_type),
    .io_grant_bits_payload_data(finisher_io_grant_bits_payload_data),
    .io_refill_ready(finisher_io_refill_ready),
    .io_refill_valid(finisher_io_refill_valid),
    .io_refill_bits_addr_beat(finisher_io_refill_bits_addr_beat),
    .io_refill_bits_client_xact_id(finisher_io_refill_bits_client_xact_id),
    .io_refill_bits_manager_xact_id(finisher_io_refill_bits_manager_xact_id),
    .io_refill_bits_is_builtin_type(finisher_io_refill_bits_is_builtin_type),
    .io_refill_bits_g_type(finisher_io_refill_bits_g_type),
    .io_refill_bits_data(finisher_io_refill_bits_data),
    .io_finish_ready(finisher_io_finish_ready),
    .io_finish_valid(finisher_io_finish_valid),
    .io_finish_bits_header_src(finisher_io_finish_bits_header_src),
    .io_finish_bits_header_dst(finisher_io_finish_bits_header_dst),
    .io_finish_bits_payload_manager_xact_id(finisher_io_finish_bits_payload_manager_xact_id),
    .io_ready(finisher_io_ready)
  );
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_network_acquire_valid = T_3339;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_probe_ready = 1'h0;
  assign io_network_release_valid = 1'h0;
  assign io_network_release_bits_header_src = GEN_1;
  assign io_network_release_bits_header_dst = GEN_2;
  assign io_network_release_bits_payload_addr_beat = GEN_3;
  assign io_network_release_bits_payload_addr_block = GEN_4;
  assign io_network_release_bits_payload_client_xact_id = GEN_5;
  assign io_network_release_bits_payload_voluntary = GEN_6;
  assign io_network_release_bits_payload_r_type = GEN_7;
  assign io_network_release_bits_payload_data = GEN_8;
  assign finisher_clk = clk;
  assign finisher_reset = reset;
  assign finisher_io_grant_valid = io_network_grant_valid;
  assign finisher_io_grant_bits_header_src = io_network_grant_bits_header_src;
  assign finisher_io_grant_bits_header_dst = io_network_grant_bits_header_dst;
  assign finisher_io_grant_bits_payload_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign finisher_io_grant_bits_payload_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign finisher_io_grant_bits_payload_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign finisher_io_grant_bits_payload_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign finisher_io_grant_bits_payload_g_type = io_network_grant_bits_payload_g_type;
  assign finisher_io_grant_bits_payload_data = io_network_grant_bits_payload_data;
  assign finisher_io_refill_ready = io_client_grant_ready;
  assign finisher_io_finish_ready = io_network_finish_ready;
  assign acq_with_header_ready = T_3340;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = 2'h1;
  assign acq_with_header_bits_header_dst = {{1'd0}, T_3338};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_3330 = GEN_0 << 6;
  assign T_3332 = 32'h80000000 <= T_3330;
  assign T_3334 = T_3330 < 32'h90000000;
  assign T_3335 = T_3332 & T_3334;
  assign T_3338 = T_3335 ? 1'h0 : 1'h1;
  assign T_3339 = acq_with_header_valid & finisher_io_ready;
  assign T_3340 = io_network_acquire_ready & finisher_io_ready;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_9[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_10[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_11[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_4 = GEN_12[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_5 = GEN_13[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_6 = GEN_14[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_7 = GEN_15[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_8 = GEN_16[63:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_9 = {1{$random}};
  GEN_10 = {1{$random}};
  GEN_11 = {1{$random}};
  GEN_12 = {1{$random}};
  GEN_13 = {1{$random}};
  GEN_14 = {1{$random}};
  GEN_15 = {1{$random}};
  GEN_16 = {2{$random}};
  end
`endif
endmodule
module ManagerTileLinkNetworkPort(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output  io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [10:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output  io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input   io_manager_grant_bits_client_xact_id,
  input  [1:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input   io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input   io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output  io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output  io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [1:0] io_network_acquire_bits_header_src,
  input  [1:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input   io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [10:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [1:0] io_network_grant_bits_header_src,
  output [1:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output  io_network_grant_bits_payload_client_xact_id,
  output [1:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [1:0] io_network_finish_bits_header_src,
  input  [1:0] io_network_finish_bits_header_dst,
  input  [1:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [1:0] io_network_probe_bits_header_src,
  output [1:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [1:0] io_network_release_bits_header_src,
  input  [1:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input   io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6043_ready;
  wire  T_6043_valid;
  wire [1:0] T_6043_bits_header_src;
  wire [1:0] T_6043_bits_header_dst;
  wire [2:0] T_6043_bits_payload_addr_beat;
  wire  T_6043_bits_payload_client_xact_id;
  wire [1:0] T_6043_bits_payload_manager_xact_id;
  wire  T_6043_bits_payload_is_builtin_type;
  wire [3:0] T_6043_bits_payload_g_type;
  wire [63:0] T_6043_bits_payload_data;
  wire  T_6043_bits_payload_client_id;
  wire  T_6598_ready;
  wire  T_6598_valid;
  wire [1:0] T_6598_bits_header_src;
  wire [1:0] T_6598_bits_header_dst;
  wire [25:0] T_6598_bits_payload_addr_block;
  wire [1:0] T_6598_bits_payload_p_type;
  wire  T_6598_bits_payload_client_id;
  wire  T_6877_ready;
  wire  T_6877_valid;
  wire [25:0] T_6877_bits_addr_block;
  wire  T_6877_bits_client_xact_id;
  wire [2:0] T_6877_bits_addr_beat;
  wire  T_6877_bits_is_builtin_type;
  wire [2:0] T_6877_bits_a_type;
  wire [10:0] T_6877_bits_union;
  wire [63:0] T_6877_bits_data;
  wire  T_6993_ready;
  wire  T_6993_valid;
  wire [2:0] T_6993_bits_addr_beat;
  wire [25:0] T_6993_bits_addr_block;
  wire  T_6993_bits_client_xact_id;
  wire  T_6993_bits_voluntary;
  wire [2:0] T_6993_bits_r_type;
  wire [63:0] T_6993_bits_data;
  wire  T_7097_ready;
  wire  T_7097_valid;
  wire [1:0] T_7097_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_6877_valid;
  assign io_manager_acquire_bits_addr_block = T_6877_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_6877_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_6877_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_6877_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_6877_bits_a_type;
  assign io_manager_acquire_bits_union = T_6877_bits_union;
  assign io_manager_acquire_bits_data = T_6877_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[0];
  assign io_manager_grant_ready = T_6043_ready;
  assign io_manager_finish_valid = T_7097_valid;
  assign io_manager_finish_bits_manager_xact_id = T_7097_bits_manager_xact_id;
  assign io_manager_probe_ready = T_6598_ready;
  assign io_manager_release_valid = T_6993_valid;
  assign io_manager_release_bits_addr_beat = T_6993_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_6993_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_6993_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_6993_bits_voluntary;
  assign io_manager_release_bits_r_type = T_6993_bits_r_type;
  assign io_manager_release_bits_data = T_6993_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[0];
  assign io_network_acquire_ready = T_6877_ready;
  assign io_network_grant_valid = T_6043_valid;
  assign io_network_grant_bits_header_src = T_6043_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6043_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6043_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6043_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6043_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6043_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6043_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6043_bits_payload_data;
  assign io_network_finish_ready = T_7097_ready;
  assign io_network_probe_valid = T_6598_valid;
  assign io_network_probe_bits_header_src = T_6598_bits_header_src;
  assign io_network_probe_bits_header_dst = T_6598_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_6598_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_6598_bits_payload_p_type;
  assign io_network_release_ready = T_6993_ready;
  assign T_6043_ready = io_network_grant_ready;
  assign T_6043_valid = io_manager_grant_valid;
  assign T_6043_bits_header_src = 2'h0;
  assign T_6043_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6043_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6043_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6043_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6043_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6043_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6043_bits_payload_data = io_manager_grant_bits_data;
  assign T_6043_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_6598_ready = io_network_probe_ready;
  assign T_6598_valid = io_manager_probe_valid;
  assign T_6598_bits_header_src = 2'h0;
  assign T_6598_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_6598_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_6598_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_6598_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_6877_ready = io_manager_acquire_ready;
  assign T_6877_valid = io_network_acquire_valid;
  assign T_6877_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_6877_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_6877_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_6877_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_6877_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_6877_bits_union = io_network_acquire_bits_payload_union;
  assign T_6877_bits_data = io_network_acquire_bits_payload_data;
  assign T_6993_ready = io_manager_release_ready;
  assign T_6993_valid = io_network_release_valid;
  assign T_6993_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_6993_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_6993_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_6993_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_6993_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_6993_bits_data = io_network_release_bits_payload_data;
  assign T_7097_ready = io_manager_finish_ready;
  assign T_7097_valid = io_network_finish_valid;
  assign T_7097_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module TileLinkEnqueuer_2(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input   io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [10:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output  io_client_grant_bits_payload_client_xact_id,
  output [1:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [1:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input   io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output  io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [10:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input   io_manager_grant_bits_payload_client_xact_id,
  input  [1:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [1:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output  io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  assign io_client_acquire_ready = io_manager_acquire_ready;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_release_ready = io_manager_release_ready;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_release_valid = io_client_release_valid;
  assign io_manager_release_bits_header_src = io_client_release_bits_header_src;
  assign io_manager_release_bits_header_dst = io_client_release_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = io_client_release_bits_payload_data;
endmodule
module ManagerTileLinkNetworkPort_1(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output  io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [10:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output  io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input   io_manager_grant_bits_client_xact_id,
  input  [1:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input   io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input   io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output  io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output  io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [1:0] io_network_acquire_bits_header_src,
  input  [1:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input   io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [10:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [1:0] io_network_grant_bits_header_src,
  output [1:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output  io_network_grant_bits_payload_client_xact_id,
  output [1:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [1:0] io_network_finish_bits_header_src,
  input  [1:0] io_network_finish_bits_header_dst,
  input  [1:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [1:0] io_network_probe_bits_header_src,
  output [1:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [1:0] io_network_release_bits_header_src,
  input  [1:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input   io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6043_ready;
  wire  T_6043_valid;
  wire [1:0] T_6043_bits_header_src;
  wire [1:0] T_6043_bits_header_dst;
  wire [2:0] T_6043_bits_payload_addr_beat;
  wire  T_6043_bits_payload_client_xact_id;
  wire [1:0] T_6043_bits_payload_manager_xact_id;
  wire  T_6043_bits_payload_is_builtin_type;
  wire [3:0] T_6043_bits_payload_g_type;
  wire [63:0] T_6043_bits_payload_data;
  wire  T_6043_bits_payload_client_id;
  wire  T_6598_ready;
  wire  T_6598_valid;
  wire [1:0] T_6598_bits_header_src;
  wire [1:0] T_6598_bits_header_dst;
  wire [25:0] T_6598_bits_payload_addr_block;
  wire [1:0] T_6598_bits_payload_p_type;
  wire  T_6598_bits_payload_client_id;
  wire  T_6877_ready;
  wire  T_6877_valid;
  wire [25:0] T_6877_bits_addr_block;
  wire  T_6877_bits_client_xact_id;
  wire [2:0] T_6877_bits_addr_beat;
  wire  T_6877_bits_is_builtin_type;
  wire [2:0] T_6877_bits_a_type;
  wire [10:0] T_6877_bits_union;
  wire [63:0] T_6877_bits_data;
  wire  T_6993_ready;
  wire  T_6993_valid;
  wire [2:0] T_6993_bits_addr_beat;
  wire [25:0] T_6993_bits_addr_block;
  wire  T_6993_bits_client_xact_id;
  wire  T_6993_bits_voluntary;
  wire [2:0] T_6993_bits_r_type;
  wire [63:0] T_6993_bits_data;
  wire  T_7097_ready;
  wire  T_7097_valid;
  wire [1:0] T_7097_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_6877_valid;
  assign io_manager_acquire_bits_addr_block = T_6877_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_6877_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_6877_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_6877_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_6877_bits_a_type;
  assign io_manager_acquire_bits_union = T_6877_bits_union;
  assign io_manager_acquire_bits_data = T_6877_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[0];
  assign io_manager_grant_ready = T_6043_ready;
  assign io_manager_finish_valid = T_7097_valid;
  assign io_manager_finish_bits_manager_xact_id = T_7097_bits_manager_xact_id;
  assign io_manager_probe_ready = T_6598_ready;
  assign io_manager_release_valid = T_6993_valid;
  assign io_manager_release_bits_addr_beat = T_6993_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_6993_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_6993_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_6993_bits_voluntary;
  assign io_manager_release_bits_r_type = T_6993_bits_r_type;
  assign io_manager_release_bits_data = T_6993_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[0];
  assign io_network_acquire_ready = T_6877_ready;
  assign io_network_grant_valid = T_6043_valid;
  assign io_network_grant_bits_header_src = T_6043_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6043_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6043_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6043_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6043_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6043_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6043_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6043_bits_payload_data;
  assign io_network_finish_ready = T_7097_ready;
  assign io_network_probe_valid = T_6598_valid;
  assign io_network_probe_bits_header_src = T_6598_bits_header_src;
  assign io_network_probe_bits_header_dst = T_6598_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_6598_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_6598_bits_payload_p_type;
  assign io_network_release_ready = T_6993_ready;
  assign T_6043_ready = io_network_grant_ready;
  assign T_6043_valid = io_manager_grant_valid;
  assign T_6043_bits_header_src = 2'h1;
  assign T_6043_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6043_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6043_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6043_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6043_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6043_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6043_bits_payload_data = io_manager_grant_bits_data;
  assign T_6043_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_6598_ready = io_network_probe_ready;
  assign T_6598_valid = io_manager_probe_valid;
  assign T_6598_bits_header_src = 2'h1;
  assign T_6598_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_6598_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_6598_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_6598_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_6877_ready = io_manager_acquire_ready;
  assign T_6877_valid = io_network_acquire_valid;
  assign T_6877_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_6877_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_6877_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_6877_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_6877_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_6877_bits_union = io_network_acquire_bits_payload_union;
  assign T_6877_bits_data = io_network_acquire_bits_payload_data;
  assign T_6993_ready = io_manager_release_ready;
  assign T_6993_valid = io_network_release_valid;
  assign T_6993_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_6993_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_6993_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_6993_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_6993_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_6993_bits_data = io_network_release_bits_payload_data;
  assign T_7097_ready = io_manager_finish_ready;
  assign T_7097_valid = io_network_finish_valid;
  assign T_7097_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module LockingRRArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input   io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [10:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input   io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [10:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input   io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [10:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input   io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [10:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output  io_out_bits_payload_client_xact_id,
  output [2:0] io_out_bits_payload_addr_beat,
  output  io_out_bits_payload_is_builtin_type,
  output [2:0] io_out_bits_payload_a_type,
  output [10:0] io_out_bits_payload_union,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire  GEN_0_bits_payload_client_xact_id;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire  GEN_0_bits_payload_is_builtin_type;
  wire [2:0] GEN_0_bits_payload_a_type;
  wire [10:0] GEN_0_bits_payload_union;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_10;
  wire  GEN_11;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [25:0] GEN_14;
  wire  GEN_15;
  wire [2:0] GEN_16;
  wire  GEN_17;
  wire [2:0] GEN_18;
  wire [10:0] GEN_19;
  wire [63:0] GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [25:0] GEN_25;
  wire  GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [2:0] GEN_29;
  wire [10:0] GEN_30;
  wire [63:0] GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire [1:0] GEN_34;
  wire [1:0] GEN_35;
  wire [25:0] GEN_36;
  wire  GEN_37;
  wire [2:0] GEN_38;
  wire  GEN_39;
  wire [2:0] GEN_40;
  wire [10:0] GEN_41;
  wire [63:0] GEN_42;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [25:0] GEN_1_bits_payload_addr_block;
  wire  GEN_1_bits_payload_client_xact_id;
  wire [2:0] GEN_1_bits_payload_addr_beat;
  wire  GEN_1_bits_payload_is_builtin_type;
  wire [2:0] GEN_1_bits_payload_a_type;
  wire [10:0] GEN_1_bits_payload_union;
  wire [63:0] GEN_1_bits_payload_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [25:0] GEN_2_bits_payload_addr_block;
  wire  GEN_2_bits_payload_client_xact_id;
  wire [2:0] GEN_2_bits_payload_addr_beat;
  wire  GEN_2_bits_payload_is_builtin_type;
  wire [2:0] GEN_2_bits_payload_a_type;
  wire [10:0] GEN_2_bits_payload_union;
  wire [63:0] GEN_2_bits_payload_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [25:0] GEN_3_bits_payload_addr_block;
  wire  GEN_3_bits_payload_client_xact_id;
  wire [2:0] GEN_3_bits_payload_addr_beat;
  wire  GEN_3_bits_payload_is_builtin_type;
  wire [2:0] GEN_3_bits_payload_a_type;
  wire [10:0] GEN_3_bits_payload_union;
  wire [63:0] GEN_3_bits_payload_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [1:0] GEN_4_bits_header_src;
  wire [1:0] GEN_4_bits_header_dst;
  wire [25:0] GEN_4_bits_payload_addr_block;
  wire  GEN_4_bits_payload_client_xact_id;
  wire [2:0] GEN_4_bits_payload_addr_beat;
  wire  GEN_4_bits_payload_is_builtin_type;
  wire [2:0] GEN_4_bits_payload_a_type;
  wire [10:0] GEN_4_bits_payload_union;
  wire [63:0] GEN_4_bits_payload_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [1:0] GEN_5_bits_header_src;
  wire [1:0] GEN_5_bits_header_dst;
  wire [25:0] GEN_5_bits_payload_addr_block;
  wire  GEN_5_bits_payload_client_xact_id;
  wire [2:0] GEN_5_bits_payload_addr_beat;
  wire  GEN_5_bits_payload_is_builtin_type;
  wire [2:0] GEN_5_bits_payload_a_type;
  wire [10:0] GEN_5_bits_payload_union;
  wire [63:0] GEN_5_bits_payload_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [1:0] GEN_6_bits_header_src;
  wire [1:0] GEN_6_bits_header_dst;
  wire [25:0] GEN_6_bits_payload_addr_block;
  wire  GEN_6_bits_payload_client_xact_id;
  wire [2:0] GEN_6_bits_payload_addr_beat;
  wire  GEN_6_bits_payload_is_builtin_type;
  wire [2:0] GEN_6_bits_payload_a_type;
  wire [10:0] GEN_6_bits_payload_union;
  wire [63:0] GEN_6_bits_payload_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [1:0] GEN_7_bits_header_src;
  wire [1:0] GEN_7_bits_header_dst;
  wire [25:0] GEN_7_bits_payload_addr_block;
  wire  GEN_7_bits_payload_client_xact_id;
  wire [2:0] GEN_7_bits_payload_addr_beat;
  wire  GEN_7_bits_payload_is_builtin_type;
  wire [2:0] GEN_7_bits_payload_a_type;
  wire [10:0] GEN_7_bits_payload_union;
  wire [63:0] GEN_7_bits_payload_data;
  wire  GEN_8_ready;
  wire  GEN_8_valid;
  wire [1:0] GEN_8_bits_header_src;
  wire [1:0] GEN_8_bits_header_dst;
  wire [25:0] GEN_8_bits_payload_addr_block;
  wire  GEN_8_bits_payload_client_xact_id;
  wire [2:0] GEN_8_bits_payload_addr_beat;
  wire  GEN_8_bits_payload_is_builtin_type;
  wire [2:0] GEN_8_bits_payload_a_type;
  wire [10:0] GEN_8_bits_payload_union;
  wire [63:0] GEN_8_bits_payload_data;
  wire  GEN_9_ready;
  wire  GEN_9_valid;
  wire [1:0] GEN_9_bits_header_src;
  wire [1:0] GEN_9_bits_header_dst;
  wire [25:0] GEN_9_bits_payload_addr_block;
  wire  GEN_9_bits_payload_client_xact_id;
  wire [2:0] GEN_9_bits_payload_addr_beat;
  wire  GEN_9_bits_payload_is_builtin_type;
  wire [2:0] GEN_9_bits_payload_a_type;
  wire [10:0] GEN_9_bits_payload_union;
  wire [63:0] GEN_9_bits_payload_data;
  reg [2:0] T_1134;
  reg [31:0] GEN_0;
  reg [1:0] T_1136;
  reg [31:0] GEN_1;
  wire  T_1138;
  wire [2:0] T_1147_0;
  wire  T_1149;
  wire  T_1150;
  wire  T_1151;
  wire  T_1152;
  wire [3:0] T_1156;
  wire [2:0] T_1157;
  wire [1:0] GEN_340;
  wire [2:0] GEN_341;
  wire [1:0] GEN_342;
  reg [1:0] lastGrant;
  reg [31:0] GEN_2;
  wire [1:0] GEN_343;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_1165;
  wire  T_1166;
  wire  T_1167;
  wire  T_1168;
  wire  T_1169;
  wire  T_1173;
  wire  T_1175;
  wire  T_1177;
  wire  T_1179;
  wire  T_1181;
  wire  T_1183;
  wire  T_1187;
  wire  T_1188;
  wire  T_1189;
  wire  T_1190;
  wire  T_1191;
  wire  T_1193;
  wire  T_1194;
  wire  T_1195;
  wire  T_1197;
  wire  T_1198;
  wire  T_1199;
  wire  T_1201;
  wire  T_1202;
  wire  T_1203;
  wire  T_1205;
  wire  T_1206;
  wire  T_1207;
  wire [1:0] GEN_344;
  wire [1:0] GEN_345;
  wire [1:0] GEN_346;
  wire [1:0] GEN_347;
  wire [1:0] GEN_348;
  wire [1:0] GEN_349;
  assign io_in_0_ready = T_1195;
  assign io_in_1_ready = T_1199;
  assign io_in_2_ready = T_1203;
  assign io_in_3_ready = T_1207;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_addr_block = GEN_3_bits_payload_addr_block;
  assign io_out_bits_payload_client_xact_id = GEN_4_bits_payload_client_xact_id;
  assign io_out_bits_payload_addr_beat = GEN_5_bits_payload_addr_beat;
  assign io_out_bits_payload_is_builtin_type = GEN_6_bits_payload_is_builtin_type;
  assign io_out_bits_payload_a_type = GEN_7_bits_payload_a_type;
  assign io_out_bits_payload_union = GEN_8_bits_payload_union;
  assign io_out_bits_payload_data = GEN_9_bits_payload_data;
  assign io_chosen = GEN_342;
  assign choice = GEN_349;
  assign GEN_0_ready = GEN_32;
  assign GEN_0_valid = GEN_33;
  assign GEN_0_bits_header_src = GEN_34;
  assign GEN_0_bits_header_dst = GEN_35;
  assign GEN_0_bits_payload_addr_block = GEN_36;
  assign GEN_0_bits_payload_client_xact_id = GEN_37;
  assign GEN_0_bits_payload_addr_beat = GEN_38;
  assign GEN_0_bits_payload_is_builtin_type = GEN_39;
  assign GEN_0_bits_payload_a_type = GEN_40;
  assign GEN_0_bits_payload_union = GEN_41;
  assign GEN_0_bits_payload_data = GEN_42;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_18 = 2'h1 == io_chosen ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign GEN_19 = 2'h1 == io_chosen ? io_in_1_bits_payload_union : io_in_0_bits_payload_union;
  assign GEN_20 = 2'h1 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_ready : GEN_10;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_valid : GEN_11;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_12;
  assign GEN_24 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_13;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_14;
  assign GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_15;
  assign GEN_27 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_16;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_17;
  assign GEN_29 = 2'h2 == io_chosen ? io_in_2_bits_payload_a_type : GEN_18;
  assign GEN_30 = 2'h2 == io_chosen ? io_in_2_bits_payload_union : GEN_19;
  assign GEN_31 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_20;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_ready : GEN_21;
  assign GEN_33 = 2'h3 == io_chosen ? io_in_3_valid : GEN_22;
  assign GEN_34 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_23;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_24;
  assign GEN_36 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_25;
  assign GEN_37 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_26;
  assign GEN_38 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_27;
  assign GEN_39 = 2'h3 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_28;
  assign GEN_40 = 2'h3 == io_chosen ? io_in_3_bits_payload_a_type : GEN_29;
  assign GEN_41 = 2'h3 == io_chosen ? io_in_3_bits_payload_union : GEN_30;
  assign GEN_42 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_31;
  assign GEN_1_ready = GEN_32;
  assign GEN_1_valid = GEN_33;
  assign GEN_1_bits_header_src = GEN_34;
  assign GEN_1_bits_header_dst = GEN_35;
  assign GEN_1_bits_payload_addr_block = GEN_36;
  assign GEN_1_bits_payload_client_xact_id = GEN_37;
  assign GEN_1_bits_payload_addr_beat = GEN_38;
  assign GEN_1_bits_payload_is_builtin_type = GEN_39;
  assign GEN_1_bits_payload_a_type = GEN_40;
  assign GEN_1_bits_payload_union = GEN_41;
  assign GEN_1_bits_payload_data = GEN_42;
  assign GEN_2_ready = GEN_32;
  assign GEN_2_valid = GEN_33;
  assign GEN_2_bits_header_src = GEN_34;
  assign GEN_2_bits_header_dst = GEN_35;
  assign GEN_2_bits_payload_addr_block = GEN_36;
  assign GEN_2_bits_payload_client_xact_id = GEN_37;
  assign GEN_2_bits_payload_addr_beat = GEN_38;
  assign GEN_2_bits_payload_is_builtin_type = GEN_39;
  assign GEN_2_bits_payload_a_type = GEN_40;
  assign GEN_2_bits_payload_union = GEN_41;
  assign GEN_2_bits_payload_data = GEN_42;
  assign GEN_3_ready = GEN_32;
  assign GEN_3_valid = GEN_33;
  assign GEN_3_bits_header_src = GEN_34;
  assign GEN_3_bits_header_dst = GEN_35;
  assign GEN_3_bits_payload_addr_block = GEN_36;
  assign GEN_3_bits_payload_client_xact_id = GEN_37;
  assign GEN_3_bits_payload_addr_beat = GEN_38;
  assign GEN_3_bits_payload_is_builtin_type = GEN_39;
  assign GEN_3_bits_payload_a_type = GEN_40;
  assign GEN_3_bits_payload_union = GEN_41;
  assign GEN_3_bits_payload_data = GEN_42;
  assign GEN_4_ready = GEN_32;
  assign GEN_4_valid = GEN_33;
  assign GEN_4_bits_header_src = GEN_34;
  assign GEN_4_bits_header_dst = GEN_35;
  assign GEN_4_bits_payload_addr_block = GEN_36;
  assign GEN_4_bits_payload_client_xact_id = GEN_37;
  assign GEN_4_bits_payload_addr_beat = GEN_38;
  assign GEN_4_bits_payload_is_builtin_type = GEN_39;
  assign GEN_4_bits_payload_a_type = GEN_40;
  assign GEN_4_bits_payload_union = GEN_41;
  assign GEN_4_bits_payload_data = GEN_42;
  assign GEN_5_ready = GEN_32;
  assign GEN_5_valid = GEN_33;
  assign GEN_5_bits_header_src = GEN_34;
  assign GEN_5_bits_header_dst = GEN_35;
  assign GEN_5_bits_payload_addr_block = GEN_36;
  assign GEN_5_bits_payload_client_xact_id = GEN_37;
  assign GEN_5_bits_payload_addr_beat = GEN_38;
  assign GEN_5_bits_payload_is_builtin_type = GEN_39;
  assign GEN_5_bits_payload_a_type = GEN_40;
  assign GEN_5_bits_payload_union = GEN_41;
  assign GEN_5_bits_payload_data = GEN_42;
  assign GEN_6_ready = GEN_32;
  assign GEN_6_valid = GEN_33;
  assign GEN_6_bits_header_src = GEN_34;
  assign GEN_6_bits_header_dst = GEN_35;
  assign GEN_6_bits_payload_addr_block = GEN_36;
  assign GEN_6_bits_payload_client_xact_id = GEN_37;
  assign GEN_6_bits_payload_addr_beat = GEN_38;
  assign GEN_6_bits_payload_is_builtin_type = GEN_39;
  assign GEN_6_bits_payload_a_type = GEN_40;
  assign GEN_6_bits_payload_union = GEN_41;
  assign GEN_6_bits_payload_data = GEN_42;
  assign GEN_7_ready = GEN_32;
  assign GEN_7_valid = GEN_33;
  assign GEN_7_bits_header_src = GEN_34;
  assign GEN_7_bits_header_dst = GEN_35;
  assign GEN_7_bits_payload_addr_block = GEN_36;
  assign GEN_7_bits_payload_client_xact_id = GEN_37;
  assign GEN_7_bits_payload_addr_beat = GEN_38;
  assign GEN_7_bits_payload_is_builtin_type = GEN_39;
  assign GEN_7_bits_payload_a_type = GEN_40;
  assign GEN_7_bits_payload_union = GEN_41;
  assign GEN_7_bits_payload_data = GEN_42;
  assign GEN_8_ready = GEN_32;
  assign GEN_8_valid = GEN_33;
  assign GEN_8_bits_header_src = GEN_34;
  assign GEN_8_bits_header_dst = GEN_35;
  assign GEN_8_bits_payload_addr_block = GEN_36;
  assign GEN_8_bits_payload_client_xact_id = GEN_37;
  assign GEN_8_bits_payload_addr_beat = GEN_38;
  assign GEN_8_bits_payload_is_builtin_type = GEN_39;
  assign GEN_8_bits_payload_a_type = GEN_40;
  assign GEN_8_bits_payload_union = GEN_41;
  assign GEN_8_bits_payload_data = GEN_42;
  assign GEN_9_ready = GEN_32;
  assign GEN_9_valid = GEN_33;
  assign GEN_9_bits_header_src = GEN_34;
  assign GEN_9_bits_header_dst = GEN_35;
  assign GEN_9_bits_payload_addr_block = GEN_36;
  assign GEN_9_bits_payload_client_xact_id = GEN_37;
  assign GEN_9_bits_payload_addr_beat = GEN_38;
  assign GEN_9_bits_payload_is_builtin_type = GEN_39;
  assign GEN_9_bits_payload_a_type = GEN_40;
  assign GEN_9_bits_payload_union = GEN_41;
  assign GEN_9_bits_payload_data = GEN_42;
  assign T_1138 = T_1134 != 3'h0;
  assign T_1147_0 = 3'h3;
  assign T_1149 = io_out_bits_payload_a_type == T_1147_0;
  assign T_1150 = io_out_bits_payload_is_builtin_type & T_1149;
  assign T_1151 = io_out_ready & io_out_valid;
  assign T_1152 = T_1151 & T_1150;
  assign T_1156 = T_1134 + 3'h1;
  assign T_1157 = T_1156[2:0];
  assign GEN_340 = T_1152 ? io_chosen : T_1136;
  assign GEN_341 = T_1152 ? T_1157 : T_1134;
  assign GEN_342 = T_1138 ? T_1136 : choice;
  assign GEN_343 = T_1151 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_1165 = validMask_1 | validMask_2;
  assign T_1166 = T_1165 | validMask_3;
  assign T_1167 = T_1166 | io_in_0_valid;
  assign T_1168 = T_1167 | io_in_1_valid;
  assign T_1169 = T_1168 | io_in_2_valid;
  assign T_1173 = validMask_1 == 1'h0;
  assign T_1175 = T_1165 == 1'h0;
  assign T_1177 = T_1166 == 1'h0;
  assign T_1179 = T_1167 == 1'h0;
  assign T_1181 = T_1168 == 1'h0;
  assign T_1183 = T_1169 == 1'h0;
  assign T_1187 = grantMask_1 | T_1179;
  assign T_1188 = T_1173 & grantMask_2;
  assign T_1189 = T_1188 | T_1181;
  assign T_1190 = T_1175 & grantMask_3;
  assign T_1191 = T_1190 | T_1183;
  assign T_1193 = T_1136 == 2'h0;
  assign T_1194 = T_1138 ? T_1193 : T_1177;
  assign T_1195 = T_1194 & io_out_ready;
  assign T_1197 = T_1136 == 2'h1;
  assign T_1198 = T_1138 ? T_1197 : T_1187;
  assign T_1199 = T_1198 & io_out_ready;
  assign T_1201 = T_1136 == 2'h2;
  assign T_1202 = T_1138 ? T_1201 : T_1189;
  assign T_1203 = T_1202 & io_out_ready;
  assign T_1205 = T_1136 == 2'h3;
  assign T_1206 = T_1138 ? T_1205 : T_1191;
  assign T_1207 = T_1206 & io_out_ready;
  assign GEN_344 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_345 = io_in_1_valid ? 2'h1 : GEN_344;
  assign GEN_346 = io_in_0_valid ? 2'h0 : GEN_345;
  assign GEN_347 = validMask_3 ? 2'h3 : GEN_346;
  assign GEN_348 = validMask_2 ? 2'h2 : GEN_347;
  assign GEN_349 = validMask_1 ? 2'h1 : GEN_348;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_1134 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_1136 = GEN_1[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1134 <= 3'h0;
    end else begin
      if(T_1152) begin
        T_1134 <= T_1157;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1152) begin
        T_1136 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1151) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input   io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [10:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input   io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [10:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input   io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [10:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input   io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [10:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output  io_out_0_bits_payload_client_xact_id,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output  io_out_0_bits_payload_is_builtin_type,
  output [2:0] io_out_0_bits_payload_a_type,
  output [10:0] io_out_0_bits_payload_union,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output  io_out_1_bits_payload_client_xact_id,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output  io_out_1_bits_payload_is_builtin_type,
  output [2:0] io_out_1_bits_payload_a_type,
  output [10:0] io_out_1_bits_payload_union,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output  io_out_2_bits_payload_client_xact_id,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output  io_out_2_bits_payload_is_builtin_type,
  output [2:0] io_out_2_bits_payload_a_type,
  output [10:0] io_out_2_bits_payload_union,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output  io_out_3_bits_payload_client_xact_id,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output  io_out_3_bits_payload_is_builtin_type,
  output [2:0] io_out_3_bits_payload_a_type,
  output [10:0] io_out_3_bits_payload_union,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire  arb_io_in_0_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_0_bits_payload_a_type;
  wire [10:0] arb_io_in_0_bits_payload_union;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire  arb_io_in_1_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_1_bits_payload_a_type;
  wire [10:0] arb_io_in_1_bits_payload_union;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire  arb_io_in_2_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_2_bits_payload_a_type;
  wire [10:0] arb_io_in_2_bits_payload_union;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire  arb_io_in_3_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_3_bits_payload_a_type;
  wire [10:0] arb_io_in_3_bits_payload_union;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire  arb_io_out_bits_payload_client_xact_id;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [2:0] arb_io_out_bits_payload_a_type;
  wire [10:0] arb_io_out_bits_payload_union;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire  GEN_0_bits_payload_client_xact_id;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire  GEN_0_bits_payload_is_builtin_type;
  wire [2:0] GEN_0_bits_payload_a_type;
  wire [10:0] GEN_0_bits_payload_union;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [25:0] GEN_5;
  wire  GEN_6;
  wire [2:0] GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [10:0] GEN_10;
  wire [63:0] GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire [25:0] GEN_16;
  wire  GEN_17;
  wire [2:0] GEN_18;
  wire  GEN_19;
  wire [2:0] GEN_20;
  wire [10:0] GEN_21;
  wire [63:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  wire [25:0] GEN_27;
  wire  GEN_28;
  wire [2:0] GEN_29;
  wire  GEN_30;
  wire [2:0] GEN_31;
  wire [10:0] GEN_32;
  wire [63:0] GEN_33;
  wire  T_1529;
  wire  T_1530;
  wire  T_1532;
  wire  T_1533;
  wire  T_1535;
  wire  T_1536;
  wire  T_1538;
  wire  T_1539;
  LockingRRArbiter arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(arb_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(arb_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(arb_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(arb_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(arb_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(arb_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(arb_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(arb_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_a_type(arb_io_out_bits_payload_a_type),
    .io_out_bits_payload_union(arb_io_out_bits_payload_union),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1530;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1533;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1536;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1539;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_3_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_a_type = io_in_0_bits_payload_a_type;
  assign arb_io_in_0_bits_payload_union = io_in_0_bits_payload_union;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_a_type = io_in_1_bits_payload_a_type;
  assign arb_io_in_1_bits_payload_union = io_in_1_bits_payload_union;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_a_type = io_in_2_bits_payload_a_type;
  assign arb_io_in_2_bits_payload_union = io_in_2_bits_payload_union;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_a_type = io_in_3_bits_payload_a_type;
  assign arb_io_in_3_bits_payload_union = io_in_3_bits_payload_union;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_23;
  assign GEN_0_valid = GEN_24;
  assign GEN_0_bits_header_src = GEN_25;
  assign GEN_0_bits_header_dst = GEN_26;
  assign GEN_0_bits_payload_addr_block = GEN_27;
  assign GEN_0_bits_payload_client_xact_id = GEN_28;
  assign GEN_0_bits_payload_addr_beat = GEN_29;
  assign GEN_0_bits_payload_is_builtin_type = GEN_30;
  assign GEN_0_bits_payload_a_type = GEN_31;
  assign GEN_0_bits_payload_union = GEN_32;
  assign GEN_0_bits_payload_data = GEN_33;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_block : io_out_0_bits_payload_addr_block;
  assign GEN_6 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_client_xact_id : io_out_0_bits_payload_client_xact_id;
  assign GEN_7 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_beat : io_out_0_bits_payload_addr_beat;
  assign GEN_8 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_is_builtin_type : io_out_0_bits_payload_is_builtin_type;
  assign GEN_9 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_a_type : io_out_0_bits_payload_a_type;
  assign GEN_10 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_union : io_out_0_bits_payload_union;
  assign GEN_11 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_data : io_out_0_bits_payload_data;
  assign GEN_12 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_13 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_14 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_15 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_16 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_block : GEN_5;
  assign GEN_17 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_client_xact_id : GEN_6;
  assign GEN_18 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_beat : GEN_7;
  assign GEN_19 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_is_builtin_type : GEN_8;
  assign GEN_20 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_a_type : GEN_9;
  assign GEN_21 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_union : GEN_10;
  assign GEN_22 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_data : GEN_11;
  assign GEN_23 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_12;
  assign GEN_24 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_13;
  assign GEN_25 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_14;
  assign GEN_26 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_15;
  assign GEN_27 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_block : GEN_16;
  assign GEN_28 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_client_xact_id : GEN_17;
  assign GEN_29 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_beat : GEN_18;
  assign GEN_30 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_is_builtin_type : GEN_19;
  assign GEN_31 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_a_type : GEN_20;
  assign GEN_32 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_union : GEN_21;
  assign GEN_33 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_data : GEN_22;
  assign T_1529 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1530 = arb_io_out_valid & T_1529;
  assign T_1532 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1533 = arb_io_out_valid & T_1532;
  assign T_1535 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1536 = arb_io_out_valid & T_1535;
  assign T_1538 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1539 = arb_io_out_valid & T_1538;
endmodule
module LockingRRArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input   io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input   io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input   io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input   io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output [25:0] io_out_bits_payload_addr_block,
  output  io_out_bits_payload_client_xact_id,
  output  io_out_bits_payload_voluntary,
  output [2:0] io_out_bits_payload_r_type,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire  GEN_0_bits_payload_client_xact_id;
  wire  GEN_0_bits_payload_voluntary;
  wire [2:0] GEN_0_bits_payload_r_type;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [2:0] GEN_13;
  wire [25:0] GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [63:0] GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  wire [2:0] GEN_23;
  wire [25:0] GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire [2:0] GEN_27;
  wire [63:0] GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire [1:0] GEN_31;
  wire [1:0] GEN_32;
  wire [2:0] GEN_33;
  wire [25:0] GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire [2:0] GEN_37;
  wire [63:0] GEN_38;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [2:0] GEN_1_bits_payload_addr_beat;
  wire [25:0] GEN_1_bits_payload_addr_block;
  wire  GEN_1_bits_payload_client_xact_id;
  wire  GEN_1_bits_payload_voluntary;
  wire [2:0] GEN_1_bits_payload_r_type;
  wire [63:0] GEN_1_bits_payload_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [2:0] GEN_2_bits_payload_addr_beat;
  wire [25:0] GEN_2_bits_payload_addr_block;
  wire  GEN_2_bits_payload_client_xact_id;
  wire  GEN_2_bits_payload_voluntary;
  wire [2:0] GEN_2_bits_payload_r_type;
  wire [63:0] GEN_2_bits_payload_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [2:0] GEN_3_bits_payload_addr_beat;
  wire [25:0] GEN_3_bits_payload_addr_block;
  wire  GEN_3_bits_payload_client_xact_id;
  wire  GEN_3_bits_payload_voluntary;
  wire [2:0] GEN_3_bits_payload_r_type;
  wire [63:0] GEN_3_bits_payload_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [1:0] GEN_4_bits_header_src;
  wire [1:0] GEN_4_bits_header_dst;
  wire [2:0] GEN_4_bits_payload_addr_beat;
  wire [25:0] GEN_4_bits_payload_addr_block;
  wire  GEN_4_bits_payload_client_xact_id;
  wire  GEN_4_bits_payload_voluntary;
  wire [2:0] GEN_4_bits_payload_r_type;
  wire [63:0] GEN_4_bits_payload_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [1:0] GEN_5_bits_header_src;
  wire [1:0] GEN_5_bits_header_dst;
  wire [2:0] GEN_5_bits_payload_addr_beat;
  wire [25:0] GEN_5_bits_payload_addr_block;
  wire  GEN_5_bits_payload_client_xact_id;
  wire  GEN_5_bits_payload_voluntary;
  wire [2:0] GEN_5_bits_payload_r_type;
  wire [63:0] GEN_5_bits_payload_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [1:0] GEN_6_bits_header_src;
  wire [1:0] GEN_6_bits_header_dst;
  wire [2:0] GEN_6_bits_payload_addr_beat;
  wire [25:0] GEN_6_bits_payload_addr_block;
  wire  GEN_6_bits_payload_client_xact_id;
  wire  GEN_6_bits_payload_voluntary;
  wire [2:0] GEN_6_bits_payload_r_type;
  wire [63:0] GEN_6_bits_payload_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [1:0] GEN_7_bits_header_src;
  wire [1:0] GEN_7_bits_header_dst;
  wire [2:0] GEN_7_bits_payload_addr_beat;
  wire [25:0] GEN_7_bits_payload_addr_block;
  wire  GEN_7_bits_payload_client_xact_id;
  wire  GEN_7_bits_payload_voluntary;
  wire [2:0] GEN_7_bits_payload_r_type;
  wire [63:0] GEN_7_bits_payload_data;
  wire  GEN_8_ready;
  wire  GEN_8_valid;
  wire [1:0] GEN_8_bits_header_src;
  wire [1:0] GEN_8_bits_header_dst;
  wire [2:0] GEN_8_bits_payload_addr_beat;
  wire [25:0] GEN_8_bits_payload_addr_block;
  wire  GEN_8_bits_payload_client_xact_id;
  wire  GEN_8_bits_payload_voluntary;
  wire [2:0] GEN_8_bits_payload_r_type;
  wire [63:0] GEN_8_bits_payload_data;
  reg [2:0] T_1100;
  reg [31:0] GEN_0;
  reg [1:0] T_1102;
  reg [31:0] GEN_1;
  wire  T_1104;
  wire  T_1106;
  wire  T_1107;
  wire  T_1108;
  wire  T_1109;
  wire  T_1110;
  wire  T_1112;
  wire  T_1113;
  wire [3:0] T_1117;
  wire [2:0] T_1118;
  wire [1:0] GEN_279;
  wire [2:0] GEN_280;
  wire [1:0] GEN_281;
  reg [1:0] lastGrant;
  reg [31:0] GEN_2;
  wire [1:0] GEN_282;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_1126;
  wire  T_1127;
  wire  T_1128;
  wire  T_1129;
  wire  T_1130;
  wire  T_1134;
  wire  T_1136;
  wire  T_1138;
  wire  T_1140;
  wire  T_1142;
  wire  T_1144;
  wire  T_1148;
  wire  T_1149;
  wire  T_1150;
  wire  T_1151;
  wire  T_1152;
  wire  T_1154;
  wire  T_1155;
  wire  T_1156;
  wire  T_1158;
  wire  T_1159;
  wire  T_1160;
  wire  T_1162;
  wire  T_1163;
  wire  T_1164;
  wire  T_1166;
  wire  T_1167;
  wire  T_1168;
  wire [1:0] GEN_283;
  wire [1:0] GEN_284;
  wire [1:0] GEN_285;
  wire [1:0] GEN_286;
  wire [1:0] GEN_287;
  wire [1:0] GEN_288;
  assign io_in_0_ready = T_1156;
  assign io_in_1_ready = T_1160;
  assign io_in_2_ready = T_1164;
  assign io_in_3_ready = T_1168;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_addr_beat = GEN_3_bits_payload_addr_beat;
  assign io_out_bits_payload_addr_block = GEN_4_bits_payload_addr_block;
  assign io_out_bits_payload_client_xact_id = GEN_5_bits_payload_client_xact_id;
  assign io_out_bits_payload_voluntary = GEN_6_bits_payload_voluntary;
  assign io_out_bits_payload_r_type = GEN_7_bits_payload_r_type;
  assign io_out_bits_payload_data = GEN_8_bits_payload_data;
  assign io_chosen = GEN_281;
  assign choice = GEN_288;
  assign GEN_0_ready = GEN_29;
  assign GEN_0_valid = GEN_30;
  assign GEN_0_bits_header_src = GEN_31;
  assign GEN_0_bits_header_dst = GEN_32;
  assign GEN_0_bits_payload_addr_beat = GEN_33;
  assign GEN_0_bits_payload_addr_block = GEN_34;
  assign GEN_0_bits_payload_client_xact_id = GEN_35;
  assign GEN_0_bits_payload_voluntary = GEN_36;
  assign GEN_0_bits_payload_r_type = GEN_37;
  assign GEN_0_bits_payload_data = GEN_38;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_payload_voluntary : io_in_0_bits_payload_voluntary;
  assign GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign GEN_18 = 2'h1 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_ready : GEN_9;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_valid : GEN_10;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_11;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_12;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_13;
  assign GEN_24 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_14;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_15;
  assign GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_payload_voluntary : GEN_16;
  assign GEN_27 = 2'h2 == io_chosen ? io_in_2_bits_payload_r_type : GEN_17;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_18;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_ready : GEN_19;
  assign GEN_30 = 2'h3 == io_chosen ? io_in_3_valid : GEN_20;
  assign GEN_31 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_21;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_22;
  assign GEN_33 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_23;
  assign GEN_34 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_24;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_25;
  assign GEN_36 = 2'h3 == io_chosen ? io_in_3_bits_payload_voluntary : GEN_26;
  assign GEN_37 = 2'h3 == io_chosen ? io_in_3_bits_payload_r_type : GEN_27;
  assign GEN_38 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_28;
  assign GEN_1_ready = GEN_29;
  assign GEN_1_valid = GEN_30;
  assign GEN_1_bits_header_src = GEN_31;
  assign GEN_1_bits_header_dst = GEN_32;
  assign GEN_1_bits_payload_addr_beat = GEN_33;
  assign GEN_1_bits_payload_addr_block = GEN_34;
  assign GEN_1_bits_payload_client_xact_id = GEN_35;
  assign GEN_1_bits_payload_voluntary = GEN_36;
  assign GEN_1_bits_payload_r_type = GEN_37;
  assign GEN_1_bits_payload_data = GEN_38;
  assign GEN_2_ready = GEN_29;
  assign GEN_2_valid = GEN_30;
  assign GEN_2_bits_header_src = GEN_31;
  assign GEN_2_bits_header_dst = GEN_32;
  assign GEN_2_bits_payload_addr_beat = GEN_33;
  assign GEN_2_bits_payload_addr_block = GEN_34;
  assign GEN_2_bits_payload_client_xact_id = GEN_35;
  assign GEN_2_bits_payload_voluntary = GEN_36;
  assign GEN_2_bits_payload_r_type = GEN_37;
  assign GEN_2_bits_payload_data = GEN_38;
  assign GEN_3_ready = GEN_29;
  assign GEN_3_valid = GEN_30;
  assign GEN_3_bits_header_src = GEN_31;
  assign GEN_3_bits_header_dst = GEN_32;
  assign GEN_3_bits_payload_addr_beat = GEN_33;
  assign GEN_3_bits_payload_addr_block = GEN_34;
  assign GEN_3_bits_payload_client_xact_id = GEN_35;
  assign GEN_3_bits_payload_voluntary = GEN_36;
  assign GEN_3_bits_payload_r_type = GEN_37;
  assign GEN_3_bits_payload_data = GEN_38;
  assign GEN_4_ready = GEN_29;
  assign GEN_4_valid = GEN_30;
  assign GEN_4_bits_header_src = GEN_31;
  assign GEN_4_bits_header_dst = GEN_32;
  assign GEN_4_bits_payload_addr_beat = GEN_33;
  assign GEN_4_bits_payload_addr_block = GEN_34;
  assign GEN_4_bits_payload_client_xact_id = GEN_35;
  assign GEN_4_bits_payload_voluntary = GEN_36;
  assign GEN_4_bits_payload_r_type = GEN_37;
  assign GEN_4_bits_payload_data = GEN_38;
  assign GEN_5_ready = GEN_29;
  assign GEN_5_valid = GEN_30;
  assign GEN_5_bits_header_src = GEN_31;
  assign GEN_5_bits_header_dst = GEN_32;
  assign GEN_5_bits_payload_addr_beat = GEN_33;
  assign GEN_5_bits_payload_addr_block = GEN_34;
  assign GEN_5_bits_payload_client_xact_id = GEN_35;
  assign GEN_5_bits_payload_voluntary = GEN_36;
  assign GEN_5_bits_payload_r_type = GEN_37;
  assign GEN_5_bits_payload_data = GEN_38;
  assign GEN_6_ready = GEN_29;
  assign GEN_6_valid = GEN_30;
  assign GEN_6_bits_header_src = GEN_31;
  assign GEN_6_bits_header_dst = GEN_32;
  assign GEN_6_bits_payload_addr_beat = GEN_33;
  assign GEN_6_bits_payload_addr_block = GEN_34;
  assign GEN_6_bits_payload_client_xact_id = GEN_35;
  assign GEN_6_bits_payload_voluntary = GEN_36;
  assign GEN_6_bits_payload_r_type = GEN_37;
  assign GEN_6_bits_payload_data = GEN_38;
  assign GEN_7_ready = GEN_29;
  assign GEN_7_valid = GEN_30;
  assign GEN_7_bits_header_src = GEN_31;
  assign GEN_7_bits_header_dst = GEN_32;
  assign GEN_7_bits_payload_addr_beat = GEN_33;
  assign GEN_7_bits_payload_addr_block = GEN_34;
  assign GEN_7_bits_payload_client_xact_id = GEN_35;
  assign GEN_7_bits_payload_voluntary = GEN_36;
  assign GEN_7_bits_payload_r_type = GEN_37;
  assign GEN_7_bits_payload_data = GEN_38;
  assign GEN_8_ready = GEN_29;
  assign GEN_8_valid = GEN_30;
  assign GEN_8_bits_header_src = GEN_31;
  assign GEN_8_bits_header_dst = GEN_32;
  assign GEN_8_bits_payload_addr_beat = GEN_33;
  assign GEN_8_bits_payload_addr_block = GEN_34;
  assign GEN_8_bits_payload_client_xact_id = GEN_35;
  assign GEN_8_bits_payload_voluntary = GEN_36;
  assign GEN_8_bits_payload_r_type = GEN_37;
  assign GEN_8_bits_payload_data = GEN_38;
  assign T_1104 = T_1100 != 3'h0;
  assign T_1106 = io_out_bits_payload_r_type == 3'h0;
  assign T_1107 = io_out_bits_payload_r_type == 3'h1;
  assign T_1108 = io_out_bits_payload_r_type == 3'h2;
  assign T_1109 = T_1106 | T_1107;
  assign T_1110 = T_1109 | T_1108;
  assign T_1112 = io_out_ready & io_out_valid;
  assign T_1113 = T_1112 & T_1110;
  assign T_1117 = T_1100 + 3'h1;
  assign T_1118 = T_1117[2:0];
  assign GEN_279 = T_1113 ? io_chosen : T_1102;
  assign GEN_280 = T_1113 ? T_1118 : T_1100;
  assign GEN_281 = T_1104 ? T_1102 : choice;
  assign GEN_282 = T_1112 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_1126 = validMask_1 | validMask_2;
  assign T_1127 = T_1126 | validMask_3;
  assign T_1128 = T_1127 | io_in_0_valid;
  assign T_1129 = T_1128 | io_in_1_valid;
  assign T_1130 = T_1129 | io_in_2_valid;
  assign T_1134 = validMask_1 == 1'h0;
  assign T_1136 = T_1126 == 1'h0;
  assign T_1138 = T_1127 == 1'h0;
  assign T_1140 = T_1128 == 1'h0;
  assign T_1142 = T_1129 == 1'h0;
  assign T_1144 = T_1130 == 1'h0;
  assign T_1148 = grantMask_1 | T_1140;
  assign T_1149 = T_1134 & grantMask_2;
  assign T_1150 = T_1149 | T_1142;
  assign T_1151 = T_1136 & grantMask_3;
  assign T_1152 = T_1151 | T_1144;
  assign T_1154 = T_1102 == 2'h0;
  assign T_1155 = T_1104 ? T_1154 : T_1138;
  assign T_1156 = T_1155 & io_out_ready;
  assign T_1158 = T_1102 == 2'h1;
  assign T_1159 = T_1104 ? T_1158 : T_1148;
  assign T_1160 = T_1159 & io_out_ready;
  assign T_1162 = T_1102 == 2'h2;
  assign T_1163 = T_1104 ? T_1162 : T_1150;
  assign T_1164 = T_1163 & io_out_ready;
  assign T_1166 = T_1102 == 2'h3;
  assign T_1167 = T_1104 ? T_1166 : T_1152;
  assign T_1168 = T_1167 & io_out_ready;
  assign GEN_283 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_284 = io_in_1_valid ? 2'h1 : GEN_283;
  assign GEN_285 = io_in_0_valid ? 2'h0 : GEN_284;
  assign GEN_286 = validMask_3 ? 2'h3 : GEN_285;
  assign GEN_287 = validMask_2 ? 2'h2 : GEN_286;
  assign GEN_288 = validMask_1 ? 2'h1 : GEN_287;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_1100 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_1102 = GEN_1[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1100 <= 3'h0;
    end else begin
      if(T_1113) begin
        T_1100 <= T_1118;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1113) begin
        T_1102 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1112) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input   io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input   io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input   io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input   io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output [25:0] io_out_0_bits_payload_addr_block,
  output  io_out_0_bits_payload_client_xact_id,
  output  io_out_0_bits_payload_voluntary,
  output [2:0] io_out_0_bits_payload_r_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output [25:0] io_out_1_bits_payload_addr_block,
  output  io_out_1_bits_payload_client_xact_id,
  output  io_out_1_bits_payload_voluntary,
  output [2:0] io_out_1_bits_payload_r_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output [25:0] io_out_2_bits_payload_addr_block,
  output  io_out_2_bits_payload_client_xact_id,
  output  io_out_2_bits_payload_voluntary,
  output [2:0] io_out_2_bits_payload_r_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output [25:0] io_out_3_bits_payload_addr_block,
  output  io_out_3_bits_payload_client_xact_id,
  output  io_out_3_bits_payload_voluntary,
  output [2:0] io_out_3_bits_payload_r_type,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire  arb_io_in_0_bits_payload_client_xact_id;
  wire  arb_io_in_0_bits_payload_voluntary;
  wire [2:0] arb_io_in_0_bits_payload_r_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire  arb_io_in_1_bits_payload_client_xact_id;
  wire  arb_io_in_1_bits_payload_voluntary;
  wire [2:0] arb_io_in_1_bits_payload_r_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire  arb_io_in_2_bits_payload_client_xact_id;
  wire  arb_io_in_2_bits_payload_voluntary;
  wire [2:0] arb_io_in_2_bits_payload_r_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire  arb_io_in_3_bits_payload_client_xact_id;
  wire  arb_io_in_3_bits_payload_voluntary;
  wire [2:0] arb_io_in_3_bits_payload_r_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire  arb_io_out_bits_payload_client_xact_id;
  wire  arb_io_out_bits_payload_voluntary;
  wire [2:0] arb_io_out_bits_payload_r_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire  GEN_0_bits_payload_client_xact_id;
  wire  GEN_0_bits_payload_voluntary;
  wire [2:0] GEN_0_bits_payload_r_type;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [2:0] GEN_5;
  wire [25:0] GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [63:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [2:0] GEN_15;
  wire [25:0] GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire [63:0] GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [2:0] GEN_25;
  wire [25:0] GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire [2:0] GEN_29;
  wire [63:0] GEN_30;
  wire  T_1483;
  wire  T_1484;
  wire  T_1486;
  wire  T_1487;
  wire  T_1489;
  wire  T_1490;
  wire  T_1492;
  wire  T_1493;
  LockingRRArbiter_1 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(arb_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(arb_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(arb_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(arb_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(arb_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(arb_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(arb_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(arb_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_voluntary(arb_io_out_bits_payload_voluntary),
    .io_out_bits_payload_r_type(arb_io_out_bits_payload_r_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1484;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_0_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1487;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_1_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1490;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_2_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1493;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_3_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_voluntary = io_in_0_bits_payload_voluntary;
  assign arb_io_in_0_bits_payload_r_type = io_in_0_bits_payload_r_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_voluntary = io_in_1_bits_payload_voluntary;
  assign arb_io_in_1_bits_payload_r_type = io_in_1_bits_payload_r_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_voluntary = io_in_2_bits_payload_voluntary;
  assign arb_io_in_2_bits_payload_r_type = io_in_2_bits_payload_r_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_voluntary = io_in_3_bits_payload_voluntary;
  assign arb_io_in_3_bits_payload_r_type = io_in_3_bits_payload_r_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_21;
  assign GEN_0_valid = GEN_22;
  assign GEN_0_bits_header_src = GEN_23;
  assign GEN_0_bits_header_dst = GEN_24;
  assign GEN_0_bits_payload_addr_beat = GEN_25;
  assign GEN_0_bits_payload_addr_block = GEN_26;
  assign GEN_0_bits_payload_client_xact_id = GEN_27;
  assign GEN_0_bits_payload_voluntary = GEN_28;
  assign GEN_0_bits_payload_r_type = GEN_29;
  assign GEN_0_bits_payload_data = GEN_30;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_beat : io_out_0_bits_payload_addr_beat;
  assign GEN_6 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_block : io_out_0_bits_payload_addr_block;
  assign GEN_7 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_client_xact_id : io_out_0_bits_payload_client_xact_id;
  assign GEN_8 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_voluntary : io_out_0_bits_payload_voluntary;
  assign GEN_9 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_r_type : io_out_0_bits_payload_r_type;
  assign GEN_10 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_data : io_out_0_bits_payload_data;
  assign GEN_11 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_12 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_13 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_14 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_15 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_beat : GEN_5;
  assign GEN_16 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_block : GEN_6;
  assign GEN_17 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_client_xact_id : GEN_7;
  assign GEN_18 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_voluntary : GEN_8;
  assign GEN_19 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_r_type : GEN_9;
  assign GEN_20 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_data : GEN_10;
  assign GEN_21 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_11;
  assign GEN_22 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_12;
  assign GEN_23 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_13;
  assign GEN_24 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_14;
  assign GEN_25 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_beat : GEN_15;
  assign GEN_26 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_block : GEN_16;
  assign GEN_27 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_client_xact_id : GEN_17;
  assign GEN_28 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_voluntary : GEN_18;
  assign GEN_29 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_r_type : GEN_19;
  assign GEN_30 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_data : GEN_20;
  assign T_1483 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1484 = arb_io_out_valid & T_1483;
  assign T_1486 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1487 = arb_io_out_valid & T_1486;
  assign T_1489 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1490 = arb_io_out_valid & T_1489;
  assign T_1492 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1493 = arb_io_out_valid & T_1492;
endmodule
module LockingRRArbiter_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_p_type,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire [1:0] GEN_0_bits_payload_p_type;
  wire  GEN_5;
  wire  GEN_6;
  wire [1:0] GEN_7;
  wire [1:0] GEN_8;
  wire [25:0] GEN_9;
  wire [1:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [25:0] GEN_15;
  wire [1:0] GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [1:0] GEN_19;
  wire [1:0] GEN_20;
  wire [25:0] GEN_21;
  wire [1:0] GEN_22;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [25:0] GEN_1_bits_payload_addr_block;
  wire [1:0] GEN_1_bits_payload_p_type;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [25:0] GEN_2_bits_payload_addr_block;
  wire [1:0] GEN_2_bits_payload_p_type;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [25:0] GEN_3_bits_payload_addr_block;
  wire [1:0] GEN_3_bits_payload_p_type;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [1:0] GEN_4_bits_header_src;
  wire [1:0] GEN_4_bits_header_dst;
  wire [25:0] GEN_4_bits_payload_addr_block;
  wire [1:0] GEN_4_bits_payload_p_type;
  wire  T_964;
  reg [1:0] lastGrant;
  reg [31:0] GEN_0;
  wire [1:0] GEN_95;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_970;
  wire  T_971;
  wire  T_972;
  wire  T_973;
  wire  T_974;
  wire  T_978;
  wire  T_980;
  wire  T_982;
  wire  T_984;
  wire  T_986;
  wire  T_988;
  wire  T_992;
  wire  T_993;
  wire  T_994;
  wire  T_995;
  wire  T_996;
  wire  T_997;
  wire  T_998;
  wire  T_999;
  wire  T_1000;
  wire [1:0] GEN_96;
  wire [1:0] GEN_97;
  wire [1:0] GEN_98;
  wire [1:0] GEN_99;
  wire [1:0] GEN_100;
  wire [1:0] GEN_101;
  assign io_in_0_ready = T_997;
  assign io_in_1_ready = T_998;
  assign io_in_2_ready = T_999;
  assign io_in_3_ready = T_1000;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_addr_block = GEN_3_bits_payload_addr_block;
  assign io_out_bits_payload_p_type = GEN_4_bits_payload_p_type;
  assign io_chosen = choice;
  assign choice = GEN_101;
  assign GEN_0_ready = GEN_17;
  assign GEN_0_valid = GEN_18;
  assign GEN_0_bits_header_src = GEN_19;
  assign GEN_0_bits_header_dst = GEN_20;
  assign GEN_0_bits_payload_addr_block = GEN_21;
  assign GEN_0_bits_payload_p_type = GEN_22;
  assign GEN_5 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_6 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_ready : GEN_5;
  assign GEN_12 = 2'h2 == io_chosen ? io_in_2_valid : GEN_6;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_7;
  assign GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_8;
  assign GEN_15 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_9;
  assign GEN_16 = 2'h2 == io_chosen ? io_in_2_bits_payload_p_type : GEN_10;
  assign GEN_17 = 2'h3 == io_chosen ? io_in_3_ready : GEN_11;
  assign GEN_18 = 2'h3 == io_chosen ? io_in_3_valid : GEN_12;
  assign GEN_19 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_13;
  assign GEN_20 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_14;
  assign GEN_21 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_15;
  assign GEN_22 = 2'h3 == io_chosen ? io_in_3_bits_payload_p_type : GEN_16;
  assign GEN_1_ready = GEN_17;
  assign GEN_1_valid = GEN_18;
  assign GEN_1_bits_header_src = GEN_19;
  assign GEN_1_bits_header_dst = GEN_20;
  assign GEN_1_bits_payload_addr_block = GEN_21;
  assign GEN_1_bits_payload_p_type = GEN_22;
  assign GEN_2_ready = GEN_17;
  assign GEN_2_valid = GEN_18;
  assign GEN_2_bits_header_src = GEN_19;
  assign GEN_2_bits_header_dst = GEN_20;
  assign GEN_2_bits_payload_addr_block = GEN_21;
  assign GEN_2_bits_payload_p_type = GEN_22;
  assign GEN_3_ready = GEN_17;
  assign GEN_3_valid = GEN_18;
  assign GEN_3_bits_header_src = GEN_19;
  assign GEN_3_bits_header_dst = GEN_20;
  assign GEN_3_bits_payload_addr_block = GEN_21;
  assign GEN_3_bits_payload_p_type = GEN_22;
  assign GEN_4_ready = GEN_17;
  assign GEN_4_valid = GEN_18;
  assign GEN_4_bits_header_src = GEN_19;
  assign GEN_4_bits_header_dst = GEN_20;
  assign GEN_4_bits_payload_addr_block = GEN_21;
  assign GEN_4_bits_payload_p_type = GEN_22;
  assign T_964 = io_out_ready & io_out_valid;
  assign GEN_95 = T_964 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_970 = validMask_1 | validMask_2;
  assign T_971 = T_970 | validMask_3;
  assign T_972 = T_971 | io_in_0_valid;
  assign T_973 = T_972 | io_in_1_valid;
  assign T_974 = T_973 | io_in_2_valid;
  assign T_978 = validMask_1 == 1'h0;
  assign T_980 = T_970 == 1'h0;
  assign T_982 = T_971 == 1'h0;
  assign T_984 = T_972 == 1'h0;
  assign T_986 = T_973 == 1'h0;
  assign T_988 = T_974 == 1'h0;
  assign T_992 = grantMask_1 | T_984;
  assign T_993 = T_978 & grantMask_2;
  assign T_994 = T_993 | T_986;
  assign T_995 = T_980 & grantMask_3;
  assign T_996 = T_995 | T_988;
  assign T_997 = T_982 & io_out_ready;
  assign T_998 = T_992 & io_out_ready;
  assign T_999 = T_994 & io_out_ready;
  assign T_1000 = T_996 & io_out_ready;
  assign GEN_96 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_97 = io_in_1_valid ? 2'h1 : GEN_96;
  assign GEN_98 = io_in_0_valid ? 2'h0 : GEN_97;
  assign GEN_99 = validMask_3 ? 2'h3 : GEN_98;
  assign GEN_100 = validMask_2 ? 2'h2 : GEN_99;
  assign GEN_101 = validMask_1 ? 2'h1 : GEN_100;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  lastGrant = GEN_0[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_964) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_p_type,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_p_type,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_p_type,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_p_type
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_p_type;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_p_type;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_p_type;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_p_type;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_p_type;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire [1:0] GEN_0_bits_payload_p_type;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [25:0] GEN_5;
  wire [1:0] GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire [1:0] GEN_9;
  wire [1:0] GEN_10;
  wire [25:0] GEN_11;
  wire [1:0] GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire [25:0] GEN_17;
  wire [1:0] GEN_18;
  wire  T_1299;
  wire  T_1300;
  wire  T_1302;
  wire  T_1303;
  wire  T_1305;
  wire  T_1306;
  wire  T_1308;
  wire  T_1309;
  LockingRRArbiter_2 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(arb_io_in_0_bits_payload_p_type),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(arb_io_in_1_bits_payload_p_type),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(arb_io_in_2_bits_payload_p_type),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(arb_io_in_3_bits_payload_p_type),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_p_type(arb_io_out_bits_payload_p_type),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1300;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_1_valid = T_1303;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_2_valid = T_1306;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_3_valid = T_1309;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_p_type = io_in_0_bits_payload_p_type;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_p_type = io_in_1_bits_payload_p_type;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_p_type = io_in_2_bits_payload_p_type;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_p_type = io_in_3_bits_payload_p_type;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_13;
  assign GEN_0_valid = GEN_14;
  assign GEN_0_bits_header_src = GEN_15;
  assign GEN_0_bits_header_dst = GEN_16;
  assign GEN_0_bits_payload_addr_block = GEN_17;
  assign GEN_0_bits_payload_p_type = GEN_18;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_block : io_out_0_bits_payload_addr_block;
  assign GEN_6 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_p_type : io_out_0_bits_payload_p_type;
  assign GEN_7 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_8 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_9 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_10 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_11 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_block : GEN_5;
  assign GEN_12 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_p_type : GEN_6;
  assign GEN_13 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_7;
  assign GEN_14 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_8;
  assign GEN_15 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_9;
  assign GEN_16 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_10;
  assign GEN_17 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_block : GEN_11;
  assign GEN_18 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_p_type : GEN_12;
  assign T_1299 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1300 = arb_io_out_valid & T_1299;
  assign T_1302 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1303 = arb_io_out_valid & T_1302;
  assign T_1305 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1306 = arb_io_out_valid & T_1305;
  assign T_1308 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1309 = arb_io_out_valid & T_1308;
endmodule
module LockingRRArbiter_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_client_xact_id,
  input  [1:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_client_xact_id,
  input  [1:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_client_xact_id,
  input  [1:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_client_xact_id,
  input  [1:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output  io_out_bits_payload_client_xact_id,
  output [1:0] io_out_bits_payload_manager_xact_id,
  output  io_out_bits_payload_is_builtin_type,
  output [3:0] io_out_bits_payload_g_type,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire  GEN_0_bits_payload_client_xact_id;
  wire [1:0] GEN_0_bits_payload_manager_xact_id;
  wire  GEN_0_bits_payload_is_builtin_type;
  wire [3:0] GEN_0_bits_payload_g_type;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [2:0] GEN_13;
  wire  GEN_14;
  wire [1:0] GEN_15;
  wire  GEN_16;
  wire [3:0] GEN_17;
  wire [63:0] GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  wire [2:0] GEN_23;
  wire  GEN_24;
  wire [1:0] GEN_25;
  wire  GEN_26;
  wire [3:0] GEN_27;
  wire [63:0] GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire [1:0] GEN_31;
  wire [1:0] GEN_32;
  wire [2:0] GEN_33;
  wire  GEN_34;
  wire [1:0] GEN_35;
  wire  GEN_36;
  wire [3:0] GEN_37;
  wire [63:0] GEN_38;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [2:0] GEN_1_bits_payload_addr_beat;
  wire  GEN_1_bits_payload_client_xact_id;
  wire [1:0] GEN_1_bits_payload_manager_xact_id;
  wire  GEN_1_bits_payload_is_builtin_type;
  wire [3:0] GEN_1_bits_payload_g_type;
  wire [63:0] GEN_1_bits_payload_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [2:0] GEN_2_bits_payload_addr_beat;
  wire  GEN_2_bits_payload_client_xact_id;
  wire [1:0] GEN_2_bits_payload_manager_xact_id;
  wire  GEN_2_bits_payload_is_builtin_type;
  wire [3:0] GEN_2_bits_payload_g_type;
  wire [63:0] GEN_2_bits_payload_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [2:0] GEN_3_bits_payload_addr_beat;
  wire  GEN_3_bits_payload_client_xact_id;
  wire [1:0] GEN_3_bits_payload_manager_xact_id;
  wire  GEN_3_bits_payload_is_builtin_type;
  wire [3:0] GEN_3_bits_payload_g_type;
  wire [63:0] GEN_3_bits_payload_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [1:0] GEN_4_bits_header_src;
  wire [1:0] GEN_4_bits_header_dst;
  wire [2:0] GEN_4_bits_payload_addr_beat;
  wire  GEN_4_bits_payload_client_xact_id;
  wire [1:0] GEN_4_bits_payload_manager_xact_id;
  wire  GEN_4_bits_payload_is_builtin_type;
  wire [3:0] GEN_4_bits_payload_g_type;
  wire [63:0] GEN_4_bits_payload_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [1:0] GEN_5_bits_header_src;
  wire [1:0] GEN_5_bits_header_dst;
  wire [2:0] GEN_5_bits_payload_addr_beat;
  wire  GEN_5_bits_payload_client_xact_id;
  wire [1:0] GEN_5_bits_payload_manager_xact_id;
  wire  GEN_5_bits_payload_is_builtin_type;
  wire [3:0] GEN_5_bits_payload_g_type;
  wire [63:0] GEN_5_bits_payload_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [1:0] GEN_6_bits_header_src;
  wire [1:0] GEN_6_bits_header_dst;
  wire [2:0] GEN_6_bits_payload_addr_beat;
  wire  GEN_6_bits_payload_client_xact_id;
  wire [1:0] GEN_6_bits_payload_manager_xact_id;
  wire  GEN_6_bits_payload_is_builtin_type;
  wire [3:0] GEN_6_bits_payload_g_type;
  wire [63:0] GEN_6_bits_payload_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [1:0] GEN_7_bits_header_src;
  wire [1:0] GEN_7_bits_header_dst;
  wire [2:0] GEN_7_bits_payload_addr_beat;
  wire  GEN_7_bits_payload_client_xact_id;
  wire [1:0] GEN_7_bits_payload_manager_xact_id;
  wire  GEN_7_bits_payload_is_builtin_type;
  wire [3:0] GEN_7_bits_payload_g_type;
  wire [63:0] GEN_7_bits_payload_data;
  wire  GEN_8_ready;
  wire  GEN_8_valid;
  wire [1:0] GEN_8_bits_header_src;
  wire [1:0] GEN_8_bits_header_dst;
  wire [2:0] GEN_8_bits_payload_addr_beat;
  wire  GEN_8_bits_payload_client_xact_id;
  wire [1:0] GEN_8_bits_payload_manager_xact_id;
  wire  GEN_8_bits_payload_is_builtin_type;
  wire [3:0] GEN_8_bits_payload_g_type;
  wire [63:0] GEN_8_bits_payload_data;
  reg [2:0] T_1100;
  reg [31:0] GEN_1;
  reg [1:0] T_1102;
  reg [31:0] GEN_2;
  wire  T_1104;
  wire [2:0] T_1112_0;
  wire [3:0] GEN_0;
  wire  T_1114;
  wire  T_1115;
  wire  T_1116;
  wire  T_1118;
  wire  T_1119;
  wire [3:0] T_1123;
  wire [2:0] T_1124;
  wire [1:0] GEN_279;
  wire [2:0] GEN_280;
  wire [1:0] GEN_281;
  reg [1:0] lastGrant;
  reg [31:0] GEN_3;
  wire [1:0] GEN_282;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_1132;
  wire  T_1133;
  wire  T_1134;
  wire  T_1135;
  wire  T_1136;
  wire  T_1140;
  wire  T_1142;
  wire  T_1144;
  wire  T_1146;
  wire  T_1148;
  wire  T_1150;
  wire  T_1154;
  wire  T_1155;
  wire  T_1156;
  wire  T_1157;
  wire  T_1158;
  wire  T_1160;
  wire  T_1161;
  wire  T_1162;
  wire  T_1164;
  wire  T_1165;
  wire  T_1166;
  wire  T_1168;
  wire  T_1169;
  wire  T_1170;
  wire  T_1172;
  wire  T_1173;
  wire  T_1174;
  wire [1:0] GEN_283;
  wire [1:0] GEN_284;
  wire [1:0] GEN_285;
  wire [1:0] GEN_286;
  wire [1:0] GEN_287;
  wire [1:0] GEN_288;
  assign io_in_0_ready = T_1162;
  assign io_in_1_ready = T_1166;
  assign io_in_2_ready = T_1170;
  assign io_in_3_ready = T_1174;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_addr_beat = GEN_3_bits_payload_addr_beat;
  assign io_out_bits_payload_client_xact_id = GEN_4_bits_payload_client_xact_id;
  assign io_out_bits_payload_manager_xact_id = GEN_5_bits_payload_manager_xact_id;
  assign io_out_bits_payload_is_builtin_type = GEN_6_bits_payload_is_builtin_type;
  assign io_out_bits_payload_g_type = GEN_7_bits_payload_g_type;
  assign io_out_bits_payload_data = GEN_8_bits_payload_data;
  assign io_chosen = GEN_281;
  assign choice = GEN_288;
  assign GEN_0_ready = GEN_29;
  assign GEN_0_valid = GEN_30;
  assign GEN_0_bits_header_src = GEN_31;
  assign GEN_0_bits_header_dst = GEN_32;
  assign GEN_0_bits_payload_addr_beat = GEN_33;
  assign GEN_0_bits_payload_client_xact_id = GEN_34;
  assign GEN_0_bits_payload_manager_xact_id = GEN_35;
  assign GEN_0_bits_payload_is_builtin_type = GEN_36;
  assign GEN_0_bits_payload_g_type = GEN_37;
  assign GEN_0_bits_payload_data = GEN_38;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign GEN_18 = 2'h1 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_ready : GEN_9;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_valid : GEN_10;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_11;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_12;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_13;
  assign GEN_24 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_14;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_15;
  assign GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_16;
  assign GEN_27 = 2'h2 == io_chosen ? io_in_2_bits_payload_g_type : GEN_17;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_18;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_ready : GEN_19;
  assign GEN_30 = 2'h3 == io_chosen ? io_in_3_valid : GEN_20;
  assign GEN_31 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_21;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_22;
  assign GEN_33 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_23;
  assign GEN_34 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_24;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_25;
  assign GEN_36 = 2'h3 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_26;
  assign GEN_37 = 2'h3 == io_chosen ? io_in_3_bits_payload_g_type : GEN_27;
  assign GEN_38 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_28;
  assign GEN_1_ready = GEN_29;
  assign GEN_1_valid = GEN_30;
  assign GEN_1_bits_header_src = GEN_31;
  assign GEN_1_bits_header_dst = GEN_32;
  assign GEN_1_bits_payload_addr_beat = GEN_33;
  assign GEN_1_bits_payload_client_xact_id = GEN_34;
  assign GEN_1_bits_payload_manager_xact_id = GEN_35;
  assign GEN_1_bits_payload_is_builtin_type = GEN_36;
  assign GEN_1_bits_payload_g_type = GEN_37;
  assign GEN_1_bits_payload_data = GEN_38;
  assign GEN_2_ready = GEN_29;
  assign GEN_2_valid = GEN_30;
  assign GEN_2_bits_header_src = GEN_31;
  assign GEN_2_bits_header_dst = GEN_32;
  assign GEN_2_bits_payload_addr_beat = GEN_33;
  assign GEN_2_bits_payload_client_xact_id = GEN_34;
  assign GEN_2_bits_payload_manager_xact_id = GEN_35;
  assign GEN_2_bits_payload_is_builtin_type = GEN_36;
  assign GEN_2_bits_payload_g_type = GEN_37;
  assign GEN_2_bits_payload_data = GEN_38;
  assign GEN_3_ready = GEN_29;
  assign GEN_3_valid = GEN_30;
  assign GEN_3_bits_header_src = GEN_31;
  assign GEN_3_bits_header_dst = GEN_32;
  assign GEN_3_bits_payload_addr_beat = GEN_33;
  assign GEN_3_bits_payload_client_xact_id = GEN_34;
  assign GEN_3_bits_payload_manager_xact_id = GEN_35;
  assign GEN_3_bits_payload_is_builtin_type = GEN_36;
  assign GEN_3_bits_payload_g_type = GEN_37;
  assign GEN_3_bits_payload_data = GEN_38;
  assign GEN_4_ready = GEN_29;
  assign GEN_4_valid = GEN_30;
  assign GEN_4_bits_header_src = GEN_31;
  assign GEN_4_bits_header_dst = GEN_32;
  assign GEN_4_bits_payload_addr_beat = GEN_33;
  assign GEN_4_bits_payload_client_xact_id = GEN_34;
  assign GEN_4_bits_payload_manager_xact_id = GEN_35;
  assign GEN_4_bits_payload_is_builtin_type = GEN_36;
  assign GEN_4_bits_payload_g_type = GEN_37;
  assign GEN_4_bits_payload_data = GEN_38;
  assign GEN_5_ready = GEN_29;
  assign GEN_5_valid = GEN_30;
  assign GEN_5_bits_header_src = GEN_31;
  assign GEN_5_bits_header_dst = GEN_32;
  assign GEN_5_bits_payload_addr_beat = GEN_33;
  assign GEN_5_bits_payload_client_xact_id = GEN_34;
  assign GEN_5_bits_payload_manager_xact_id = GEN_35;
  assign GEN_5_bits_payload_is_builtin_type = GEN_36;
  assign GEN_5_bits_payload_g_type = GEN_37;
  assign GEN_5_bits_payload_data = GEN_38;
  assign GEN_6_ready = GEN_29;
  assign GEN_6_valid = GEN_30;
  assign GEN_6_bits_header_src = GEN_31;
  assign GEN_6_bits_header_dst = GEN_32;
  assign GEN_6_bits_payload_addr_beat = GEN_33;
  assign GEN_6_bits_payload_client_xact_id = GEN_34;
  assign GEN_6_bits_payload_manager_xact_id = GEN_35;
  assign GEN_6_bits_payload_is_builtin_type = GEN_36;
  assign GEN_6_bits_payload_g_type = GEN_37;
  assign GEN_6_bits_payload_data = GEN_38;
  assign GEN_7_ready = GEN_29;
  assign GEN_7_valid = GEN_30;
  assign GEN_7_bits_header_src = GEN_31;
  assign GEN_7_bits_header_dst = GEN_32;
  assign GEN_7_bits_payload_addr_beat = GEN_33;
  assign GEN_7_bits_payload_client_xact_id = GEN_34;
  assign GEN_7_bits_payload_manager_xact_id = GEN_35;
  assign GEN_7_bits_payload_is_builtin_type = GEN_36;
  assign GEN_7_bits_payload_g_type = GEN_37;
  assign GEN_7_bits_payload_data = GEN_38;
  assign GEN_8_ready = GEN_29;
  assign GEN_8_valid = GEN_30;
  assign GEN_8_bits_header_src = GEN_31;
  assign GEN_8_bits_header_dst = GEN_32;
  assign GEN_8_bits_payload_addr_beat = GEN_33;
  assign GEN_8_bits_payload_client_xact_id = GEN_34;
  assign GEN_8_bits_payload_manager_xact_id = GEN_35;
  assign GEN_8_bits_payload_is_builtin_type = GEN_36;
  assign GEN_8_bits_payload_g_type = GEN_37;
  assign GEN_8_bits_payload_data = GEN_38;
  assign T_1104 = T_1100 != 3'h0;
  assign T_1112_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_1112_0};
  assign T_1114 = io_out_bits_payload_g_type == GEN_0;
  assign T_1115 = io_out_bits_payload_g_type == 4'h0;
  assign T_1116 = io_out_bits_payload_is_builtin_type ? T_1114 : T_1115;
  assign T_1118 = io_out_ready & io_out_valid;
  assign T_1119 = T_1118 & T_1116;
  assign T_1123 = T_1100 + 3'h1;
  assign T_1124 = T_1123[2:0];
  assign GEN_279 = T_1119 ? io_chosen : T_1102;
  assign GEN_280 = T_1119 ? T_1124 : T_1100;
  assign GEN_281 = T_1104 ? T_1102 : choice;
  assign GEN_282 = T_1118 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_1132 = validMask_1 | validMask_2;
  assign T_1133 = T_1132 | validMask_3;
  assign T_1134 = T_1133 | io_in_0_valid;
  assign T_1135 = T_1134 | io_in_1_valid;
  assign T_1136 = T_1135 | io_in_2_valid;
  assign T_1140 = validMask_1 == 1'h0;
  assign T_1142 = T_1132 == 1'h0;
  assign T_1144 = T_1133 == 1'h0;
  assign T_1146 = T_1134 == 1'h0;
  assign T_1148 = T_1135 == 1'h0;
  assign T_1150 = T_1136 == 1'h0;
  assign T_1154 = grantMask_1 | T_1146;
  assign T_1155 = T_1140 & grantMask_2;
  assign T_1156 = T_1155 | T_1148;
  assign T_1157 = T_1142 & grantMask_3;
  assign T_1158 = T_1157 | T_1150;
  assign T_1160 = T_1102 == 2'h0;
  assign T_1161 = T_1104 ? T_1160 : T_1144;
  assign T_1162 = T_1161 & io_out_ready;
  assign T_1164 = T_1102 == 2'h1;
  assign T_1165 = T_1104 ? T_1164 : T_1154;
  assign T_1166 = T_1165 & io_out_ready;
  assign T_1168 = T_1102 == 2'h2;
  assign T_1169 = T_1104 ? T_1168 : T_1156;
  assign T_1170 = T_1169 & io_out_ready;
  assign T_1172 = T_1102 == 2'h3;
  assign T_1173 = T_1104 ? T_1172 : T_1158;
  assign T_1174 = T_1173 & io_out_ready;
  assign GEN_283 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_284 = io_in_1_valid ? 2'h1 : GEN_283;
  assign GEN_285 = io_in_0_valid ? 2'h0 : GEN_284;
  assign GEN_286 = validMask_3 ? 2'h3 : GEN_285;
  assign GEN_287 = validMask_2 ? 2'h2 : GEN_286;
  assign GEN_288 = validMask_1 ? 2'h1 : GEN_287;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_1100 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_1102 = GEN_2[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  lastGrant = GEN_3[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1100 <= 3'h0;
    end else begin
      if(T_1119) begin
        T_1100 <= T_1124;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1119) begin
        T_1102 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1118) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_client_xact_id,
  input  [1:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_client_xact_id,
  input  [1:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_client_xact_id,
  input  [1:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_client_xact_id,
  input  [1:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output  io_out_0_bits_payload_client_xact_id,
  output [1:0] io_out_0_bits_payload_manager_xact_id,
  output  io_out_0_bits_payload_is_builtin_type,
  output [3:0] io_out_0_bits_payload_g_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output  io_out_1_bits_payload_client_xact_id,
  output [1:0] io_out_1_bits_payload_manager_xact_id,
  output  io_out_1_bits_payload_is_builtin_type,
  output [3:0] io_out_1_bits_payload_g_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output  io_out_2_bits_payload_client_xact_id,
  output [1:0] io_out_2_bits_payload_manager_xact_id,
  output  io_out_2_bits_payload_is_builtin_type,
  output [3:0] io_out_2_bits_payload_g_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output  io_out_3_bits_payload_client_xact_id,
  output [1:0] io_out_3_bits_payload_manager_xact_id,
  output  io_out_3_bits_payload_is_builtin_type,
  output [3:0] io_out_3_bits_payload_g_type,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire  arb_io_in_0_bits_payload_client_xact_id;
  wire [1:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_0_bits_payload_g_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire  arb_io_in_1_bits_payload_client_xact_id;
  wire [1:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_1_bits_payload_g_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire  arb_io_in_2_bits_payload_client_xact_id;
  wire [1:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_2_bits_payload_g_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire  arb_io_in_3_bits_payload_client_xact_id;
  wire [1:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_3_bits_payload_g_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire  arb_io_out_bits_payload_client_xact_id;
  wire [1:0] arb_io_out_bits_payload_manager_xact_id;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [3:0] arb_io_out_bits_payload_g_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire  GEN_0_bits_payload_client_xact_id;
  wire [1:0] GEN_0_bits_payload_manager_xact_id;
  wire  GEN_0_bits_payload_is_builtin_type;
  wire [3:0] GEN_0_bits_payload_g_type;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [2:0] GEN_5;
  wire  GEN_6;
  wire [1:0] GEN_7;
  wire  GEN_8;
  wire [3:0] GEN_9;
  wire [63:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  wire [1:0] GEN_17;
  wire  GEN_18;
  wire [3:0] GEN_19;
  wire [63:0] GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [2:0] GEN_25;
  wire  GEN_26;
  wire [1:0] GEN_27;
  wire  GEN_28;
  wire [3:0] GEN_29;
  wire [63:0] GEN_30;
  wire  T_1483;
  wire  T_1484;
  wire  T_1486;
  wire  T_1487;
  wire  T_1489;
  wire  T_1490;
  wire  T_1492;
  wire  T_1493;
  LockingRRArbiter_3 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(arb_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(arb_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(arb_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(arb_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_g_type(arb_io_out_bits_payload_g_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1484;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1487;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1490;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1493;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_g_type = io_in_0_bits_payload_g_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_g_type = io_in_1_bits_payload_g_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_g_type = io_in_2_bits_payload_g_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_g_type = io_in_3_bits_payload_g_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_21;
  assign GEN_0_valid = GEN_22;
  assign GEN_0_bits_header_src = GEN_23;
  assign GEN_0_bits_header_dst = GEN_24;
  assign GEN_0_bits_payload_addr_beat = GEN_25;
  assign GEN_0_bits_payload_client_xact_id = GEN_26;
  assign GEN_0_bits_payload_manager_xact_id = GEN_27;
  assign GEN_0_bits_payload_is_builtin_type = GEN_28;
  assign GEN_0_bits_payload_g_type = GEN_29;
  assign GEN_0_bits_payload_data = GEN_30;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_beat : io_out_0_bits_payload_addr_beat;
  assign GEN_6 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_client_xact_id : io_out_0_bits_payload_client_xact_id;
  assign GEN_7 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_manager_xact_id : io_out_0_bits_payload_manager_xact_id;
  assign GEN_8 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_is_builtin_type : io_out_0_bits_payload_is_builtin_type;
  assign GEN_9 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_g_type : io_out_0_bits_payload_g_type;
  assign GEN_10 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_data : io_out_0_bits_payload_data;
  assign GEN_11 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_12 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_13 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_14 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_15 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_beat : GEN_5;
  assign GEN_16 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_client_xact_id : GEN_6;
  assign GEN_17 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_manager_xact_id : GEN_7;
  assign GEN_18 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_is_builtin_type : GEN_8;
  assign GEN_19 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_g_type : GEN_9;
  assign GEN_20 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_data : GEN_10;
  assign GEN_21 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_11;
  assign GEN_22 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_12;
  assign GEN_23 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_13;
  assign GEN_24 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_14;
  assign GEN_25 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_beat : GEN_15;
  assign GEN_26 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_client_xact_id : GEN_16;
  assign GEN_27 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_manager_xact_id : GEN_17;
  assign GEN_28 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_is_builtin_type : GEN_18;
  assign GEN_29 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_g_type : GEN_19;
  assign GEN_30 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_data : GEN_20;
  assign T_1483 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1484 = arb_io_out_valid & T_1483;
  assign T_1486 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1487 = arb_io_out_valid & T_1486;
  assign T_1489 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1490 = arb_io_out_valid & T_1489;
  assign T_1492 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1493 = arb_io_out_valid & T_1492;
endmodule
module LockingRRArbiter_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [1:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [1:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [1:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [1:0] io_in_3_bits_payload_manager_xact_id,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [1:0] io_out_bits_payload_manager_xact_id,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [1:0] GEN_0_bits_payload_manager_xact_id;
  wire  GEN_4;
  wire  GEN_5;
  wire [1:0] GEN_6;
  wire [1:0] GEN_7;
  wire [1:0] GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [1:0] GEN_1_bits_payload_manager_xact_id;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [1:0] GEN_2_bits_payload_manager_xact_id;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [1:0] GEN_3_bits_payload_manager_xact_id;
  wire  T_930;
  reg [1:0] lastGrant;
  reg [31:0] GEN_0;
  wire [1:0] GEN_64;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_936;
  wire  T_937;
  wire  T_938;
  wire  T_939;
  wire  T_940;
  wire  T_944;
  wire  T_946;
  wire  T_948;
  wire  T_950;
  wire  T_952;
  wire  T_954;
  wire  T_958;
  wire  T_959;
  wire  T_960;
  wire  T_961;
  wire  T_962;
  wire  T_963;
  wire  T_964;
  wire  T_965;
  wire  T_966;
  wire [1:0] GEN_65;
  wire [1:0] GEN_66;
  wire [1:0] GEN_67;
  wire [1:0] GEN_68;
  wire [1:0] GEN_69;
  wire [1:0] GEN_70;
  assign io_in_0_ready = T_963;
  assign io_in_1_ready = T_964;
  assign io_in_2_ready = T_965;
  assign io_in_3_ready = T_966;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_manager_xact_id = GEN_3_bits_payload_manager_xact_id;
  assign io_chosen = choice;
  assign choice = GEN_70;
  assign GEN_0_ready = GEN_14;
  assign GEN_0_valid = GEN_15;
  assign GEN_0_bits_header_src = GEN_16;
  assign GEN_0_bits_header_dst = GEN_17;
  assign GEN_0_bits_payload_manager_xact_id = GEN_18;
  assign GEN_4 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_5 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_6 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_9 = 2'h2 == io_chosen ? io_in_2_ready : GEN_4;
  assign GEN_10 = 2'h2 == io_chosen ? io_in_2_valid : GEN_5;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_6;
  assign GEN_12 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_7;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_8;
  assign GEN_14 = 2'h3 == io_chosen ? io_in_3_ready : GEN_9;
  assign GEN_15 = 2'h3 == io_chosen ? io_in_3_valid : GEN_10;
  assign GEN_16 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_11;
  assign GEN_17 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_12;
  assign GEN_18 = 2'h3 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_13;
  assign GEN_1_ready = GEN_14;
  assign GEN_1_valid = GEN_15;
  assign GEN_1_bits_header_src = GEN_16;
  assign GEN_1_bits_header_dst = GEN_17;
  assign GEN_1_bits_payload_manager_xact_id = GEN_18;
  assign GEN_2_ready = GEN_14;
  assign GEN_2_valid = GEN_15;
  assign GEN_2_bits_header_src = GEN_16;
  assign GEN_2_bits_header_dst = GEN_17;
  assign GEN_2_bits_payload_manager_xact_id = GEN_18;
  assign GEN_3_ready = GEN_14;
  assign GEN_3_valid = GEN_15;
  assign GEN_3_bits_header_src = GEN_16;
  assign GEN_3_bits_header_dst = GEN_17;
  assign GEN_3_bits_payload_manager_xact_id = GEN_18;
  assign T_930 = io_out_ready & io_out_valid;
  assign GEN_64 = T_930 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_936 = validMask_1 | validMask_2;
  assign T_937 = T_936 | validMask_3;
  assign T_938 = T_937 | io_in_0_valid;
  assign T_939 = T_938 | io_in_1_valid;
  assign T_940 = T_939 | io_in_2_valid;
  assign T_944 = validMask_1 == 1'h0;
  assign T_946 = T_936 == 1'h0;
  assign T_948 = T_937 == 1'h0;
  assign T_950 = T_938 == 1'h0;
  assign T_952 = T_939 == 1'h0;
  assign T_954 = T_940 == 1'h0;
  assign T_958 = grantMask_1 | T_950;
  assign T_959 = T_944 & grantMask_2;
  assign T_960 = T_959 | T_952;
  assign T_961 = T_946 & grantMask_3;
  assign T_962 = T_961 | T_954;
  assign T_963 = T_948 & io_out_ready;
  assign T_964 = T_958 & io_out_ready;
  assign T_965 = T_960 & io_out_ready;
  assign T_966 = T_962 & io_out_ready;
  assign GEN_65 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_66 = io_in_1_valid ? 2'h1 : GEN_65;
  assign GEN_67 = io_in_0_valid ? 2'h0 : GEN_66;
  assign GEN_68 = validMask_3 ? 2'h3 : GEN_67;
  assign GEN_69 = validMask_2 ? 2'h2 : GEN_68;
  assign GEN_70 = validMask_1 ? 2'h1 : GEN_69;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  lastGrant = GEN_0[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_930) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [1:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [1:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [1:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [1:0] io_in_3_bits_payload_manager_xact_id,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [1:0] io_out_0_bits_payload_manager_xact_id,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [1:0] io_out_1_bits_payload_manager_xact_id,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [1:0] io_out_2_bits_payload_manager_xact_id,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [1:0] io_out_3_bits_payload_manager_xact_id
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [1:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [1:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [1:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [1:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [1:0] arb_io_out_bits_payload_manager_xact_id;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [1:0] GEN_0_bits_payload_manager_xact_id;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [1:0] GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [1:0] GEN_8;
  wire [1:0] GEN_9;
  wire [1:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire  T_1253;
  wire  T_1254;
  wire  T_1256;
  wire  T_1257;
  wire  T_1259;
  wire  T_1260;
  wire  T_1262;
  wire  T_1263;
  LockingRRArbiter_4 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1254;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_valid = T_1257;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_valid = T_1260;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_valid = T_1263;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_11;
  assign GEN_0_valid = GEN_12;
  assign GEN_0_bits_header_src = GEN_13;
  assign GEN_0_bits_header_dst = GEN_14;
  assign GEN_0_bits_payload_manager_xact_id = GEN_15;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_manager_xact_id : io_out_0_bits_payload_manager_xact_id;
  assign GEN_6 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_7 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_8 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_9 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_10 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_manager_xact_id : GEN_5;
  assign GEN_11 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_6;
  assign GEN_12 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_7;
  assign GEN_13 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_8;
  assign GEN_14 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_9;
  assign GEN_15 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_manager_xact_id : GEN_10;
  assign T_1253 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1254 = arb_io_out_valid & T_1253;
  assign T_1256 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1257 = arb_io_out_valid & T_1256;
  assign T_1259 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1260 = arb_io_out_valid & T_1259;
  assign T_1262 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1263 = arb_io_out_valid & T_1262;
endmodule
module PortedTileLinkCrossbar(
  input   clk,
  input   reset,
  output  io_clients_cached_0_acquire_ready,
  input   io_clients_cached_0_acquire_valid,
  input  [25:0] io_clients_cached_0_acquire_bits_addr_block,
  input   io_clients_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_cached_0_acquire_bits_addr_beat,
  input   io_clients_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_cached_0_acquire_bits_a_type,
  input  [10:0] io_clients_cached_0_acquire_bits_union,
  input  [63:0] io_clients_cached_0_acquire_bits_data,
  input   io_clients_cached_0_probe_ready,
  output  io_clients_cached_0_probe_valid,
  output [25:0] io_clients_cached_0_probe_bits_addr_block,
  output [1:0] io_clients_cached_0_probe_bits_p_type,
  output  io_clients_cached_0_release_ready,
  input   io_clients_cached_0_release_valid,
  input  [2:0] io_clients_cached_0_release_bits_addr_beat,
  input  [25:0] io_clients_cached_0_release_bits_addr_block,
  input   io_clients_cached_0_release_bits_client_xact_id,
  input   io_clients_cached_0_release_bits_voluntary,
  input  [2:0] io_clients_cached_0_release_bits_r_type,
  input  [63:0] io_clients_cached_0_release_bits_data,
  input   io_clients_cached_0_grant_ready,
  output  io_clients_cached_0_grant_valid,
  output [2:0] io_clients_cached_0_grant_bits_addr_beat,
  output  io_clients_cached_0_grant_bits_client_xact_id,
  output [1:0] io_clients_cached_0_grant_bits_manager_xact_id,
  output  io_clients_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_cached_0_grant_bits_g_type,
  output [63:0] io_clients_cached_0_grant_bits_data,
  output  io_clients_cached_0_grant_bits_manager_id,
  output  io_clients_cached_0_finish_ready,
  input   io_clients_cached_0_finish_valid,
  input  [1:0] io_clients_cached_0_finish_bits_manager_xact_id,
  input   io_clients_cached_0_finish_bits_manager_id,
  output  io_clients_uncached_0_acquire_ready,
  input   io_clients_uncached_0_acquire_valid,
  input  [25:0] io_clients_uncached_0_acquire_bits_addr_block,
  input   io_clients_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_uncached_0_acquire_bits_addr_beat,
  input   io_clients_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_uncached_0_acquire_bits_a_type,
  input  [10:0] io_clients_uncached_0_acquire_bits_union,
  input  [63:0] io_clients_uncached_0_acquire_bits_data,
  input   io_clients_uncached_0_grant_ready,
  output  io_clients_uncached_0_grant_valid,
  output [2:0] io_clients_uncached_0_grant_bits_addr_beat,
  output  io_clients_uncached_0_grant_bits_client_xact_id,
  output [1:0] io_clients_uncached_0_grant_bits_manager_xact_id,
  output  io_clients_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_uncached_0_grant_bits_g_type,
  output [63:0] io_clients_uncached_0_grant_bits_data,
  input   io_managers_0_acquire_ready,
  output  io_managers_0_acquire_valid,
  output [25:0] io_managers_0_acquire_bits_addr_block,
  output  io_managers_0_acquire_bits_client_xact_id,
  output [2:0] io_managers_0_acquire_bits_addr_beat,
  output  io_managers_0_acquire_bits_is_builtin_type,
  output [2:0] io_managers_0_acquire_bits_a_type,
  output [10:0] io_managers_0_acquire_bits_union,
  output [63:0] io_managers_0_acquire_bits_data,
  output  io_managers_0_acquire_bits_client_id,
  output  io_managers_0_grant_ready,
  input   io_managers_0_grant_valid,
  input  [2:0] io_managers_0_grant_bits_addr_beat,
  input   io_managers_0_grant_bits_client_xact_id,
  input  [1:0] io_managers_0_grant_bits_manager_xact_id,
  input   io_managers_0_grant_bits_is_builtin_type,
  input  [3:0] io_managers_0_grant_bits_g_type,
  input  [63:0] io_managers_0_grant_bits_data,
  input   io_managers_0_grant_bits_client_id,
  input   io_managers_0_finish_ready,
  output  io_managers_0_finish_valid,
  output [1:0] io_managers_0_finish_bits_manager_xact_id,
  output  io_managers_0_probe_ready,
  input   io_managers_0_probe_valid,
  input  [25:0] io_managers_0_probe_bits_addr_block,
  input  [1:0] io_managers_0_probe_bits_p_type,
  input   io_managers_0_probe_bits_client_id,
  input   io_managers_0_release_ready,
  output  io_managers_0_release_valid,
  output [2:0] io_managers_0_release_bits_addr_beat,
  output [25:0] io_managers_0_release_bits_addr_block,
  output  io_managers_0_release_bits_client_xact_id,
  output  io_managers_0_release_bits_voluntary,
  output [2:0] io_managers_0_release_bits_r_type,
  output [63:0] io_managers_0_release_bits_data,
  output  io_managers_0_release_bits_client_id,
  input   io_managers_1_acquire_ready,
  output  io_managers_1_acquire_valid,
  output [25:0] io_managers_1_acquire_bits_addr_block,
  output  io_managers_1_acquire_bits_client_xact_id,
  output [2:0] io_managers_1_acquire_bits_addr_beat,
  output  io_managers_1_acquire_bits_is_builtin_type,
  output [2:0] io_managers_1_acquire_bits_a_type,
  output [10:0] io_managers_1_acquire_bits_union,
  output [63:0] io_managers_1_acquire_bits_data,
  output  io_managers_1_acquire_bits_client_id,
  output  io_managers_1_grant_ready,
  input   io_managers_1_grant_valid,
  input  [2:0] io_managers_1_grant_bits_addr_beat,
  input   io_managers_1_grant_bits_client_xact_id,
  input  [1:0] io_managers_1_grant_bits_manager_xact_id,
  input   io_managers_1_grant_bits_is_builtin_type,
  input  [3:0] io_managers_1_grant_bits_g_type,
  input  [63:0] io_managers_1_grant_bits_data,
  input   io_managers_1_grant_bits_client_id,
  input   io_managers_1_finish_ready,
  output  io_managers_1_finish_valid,
  output [1:0] io_managers_1_finish_bits_manager_xact_id,
  output  io_managers_1_probe_ready,
  input   io_managers_1_probe_valid,
  input  [25:0] io_managers_1_probe_bits_addr_block,
  input  [1:0] io_managers_1_probe_bits_p_type,
  input   io_managers_1_probe_bits_client_id,
  input   io_managers_1_release_ready,
  output  io_managers_1_release_valid,
  output [2:0] io_managers_1_release_bits_addr_beat,
  output [25:0] io_managers_1_release_bits_addr_block,
  output  io_managers_1_release_bits_client_xact_id,
  output  io_managers_1_release_bits_voluntary,
  output [2:0] io_managers_1_release_bits_r_type,
  output [63:0] io_managers_1_release_bits_data,
  output  io_managers_1_release_bits_client_id
);
  wire  TileLinkEnqueuer_4_clk;
  wire  TileLinkEnqueuer_4_reset;
  wire  TileLinkEnqueuer_4_io_client_acquire_ready;
  wire  TileLinkEnqueuer_4_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_client_grant_ready;
  wire  TileLinkEnqueuer_4_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_client_finish_ready;
  wire  TileLinkEnqueuer_4_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_client_probe_ready;
  wire  TileLinkEnqueuer_4_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_io_client_release_ready;
  wire  TileLinkEnqueuer_4_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_4_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_grant_ready;
  wire  TileLinkEnqueuer_4_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_finish_ready;
  wire  TileLinkEnqueuer_4_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_probe_ready;
  wire  TileLinkEnqueuer_4_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_io_manager_release_ready;
  wire  TileLinkEnqueuer_4_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_clk;
  wire  ClientTileLinkNetworkPort_1_reset;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_valid;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type;
  wire [10:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_union;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_probe_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_probe_valid;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  wire  ClientTileLinkNetworkPort_1_io_client_release_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_release_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block;
  wire  ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_release_bits_r_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_release_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire [10:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_io_network_finish_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_finish_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_probe_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_probe_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type;
  wire  ClientTileLinkNetworkPort_1_io_network_release_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_release_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire  ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_clk;
  wire  TileLinkEnqueuer_1_1_reset;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_1_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_1_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_1_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_1_1_io_client_release_ready;
  wire  TileLinkEnqueuer_1_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_1_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_clk;
  wire  ClientUncachedTileLinkNetworkPort_1_reset;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire [10:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_clk;
  wire  ManagerTileLinkNetworkPort_2_reset;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type;
  wire [10:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type;
  wire [10:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_probe_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_clk;
  wire  TileLinkEnqueuer_2_1_reset;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_2_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_2_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_2_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_2_1_io_client_release_ready;
  wire  TileLinkEnqueuer_2_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_2_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_clk;
  wire  ManagerTileLinkNetworkPort_1_1_reset;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type;
  wire [10:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type;
  wire [10:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_probe_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_clk;
  wire  TileLinkEnqueuer_3_1_reset;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_3_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_3_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_3_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_3_1_io_client_release_ready;
  wire  TileLinkEnqueuer_3_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_3_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data;
  wire  acqNet_clk;
  wire  acqNet_reset;
  wire  acqNet_io_in_0_ready;
  wire  acqNet_io_in_0_valid;
  wire [1:0] acqNet_io_in_0_bits_header_src;
  wire [1:0] acqNet_io_in_0_bits_header_dst;
  wire [25:0] acqNet_io_in_0_bits_payload_addr_block;
  wire  acqNet_io_in_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_0_bits_payload_addr_beat;
  wire  acqNet_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_0_bits_payload_a_type;
  wire [10:0] acqNet_io_in_0_bits_payload_union;
  wire [63:0] acqNet_io_in_0_bits_payload_data;
  wire  acqNet_io_in_1_ready;
  wire  acqNet_io_in_1_valid;
  wire [1:0] acqNet_io_in_1_bits_header_src;
  wire [1:0] acqNet_io_in_1_bits_header_dst;
  wire [25:0] acqNet_io_in_1_bits_payload_addr_block;
  wire  acqNet_io_in_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_1_bits_payload_addr_beat;
  wire  acqNet_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_1_bits_payload_a_type;
  wire [10:0] acqNet_io_in_1_bits_payload_union;
  wire [63:0] acqNet_io_in_1_bits_payload_data;
  wire  acqNet_io_in_2_ready;
  wire  acqNet_io_in_2_valid;
  wire [1:0] acqNet_io_in_2_bits_header_src;
  wire [1:0] acqNet_io_in_2_bits_header_dst;
  wire [25:0] acqNet_io_in_2_bits_payload_addr_block;
  wire  acqNet_io_in_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_2_bits_payload_addr_beat;
  wire  acqNet_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_2_bits_payload_a_type;
  wire [10:0] acqNet_io_in_2_bits_payload_union;
  wire [63:0] acqNet_io_in_2_bits_payload_data;
  wire  acqNet_io_in_3_ready;
  wire  acqNet_io_in_3_valid;
  wire [1:0] acqNet_io_in_3_bits_header_src;
  wire [1:0] acqNet_io_in_3_bits_header_dst;
  wire [25:0] acqNet_io_in_3_bits_payload_addr_block;
  wire  acqNet_io_in_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_3_bits_payload_addr_beat;
  wire  acqNet_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_3_bits_payload_a_type;
  wire [10:0] acqNet_io_in_3_bits_payload_union;
  wire [63:0] acqNet_io_in_3_bits_payload_data;
  wire  acqNet_io_out_0_ready;
  wire  acqNet_io_out_0_valid;
  wire [1:0] acqNet_io_out_0_bits_header_src;
  wire [1:0] acqNet_io_out_0_bits_header_dst;
  wire [25:0] acqNet_io_out_0_bits_payload_addr_block;
  wire  acqNet_io_out_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_0_bits_payload_addr_beat;
  wire  acqNet_io_out_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_0_bits_payload_a_type;
  wire [10:0] acqNet_io_out_0_bits_payload_union;
  wire [63:0] acqNet_io_out_0_bits_payload_data;
  wire  acqNet_io_out_1_ready;
  wire  acqNet_io_out_1_valid;
  wire [1:0] acqNet_io_out_1_bits_header_src;
  wire [1:0] acqNet_io_out_1_bits_header_dst;
  wire [25:0] acqNet_io_out_1_bits_payload_addr_block;
  wire  acqNet_io_out_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_1_bits_payload_addr_beat;
  wire  acqNet_io_out_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_1_bits_payload_a_type;
  wire [10:0] acqNet_io_out_1_bits_payload_union;
  wire [63:0] acqNet_io_out_1_bits_payload_data;
  wire  acqNet_io_out_2_ready;
  wire  acqNet_io_out_2_valid;
  wire [1:0] acqNet_io_out_2_bits_header_src;
  wire [1:0] acqNet_io_out_2_bits_header_dst;
  wire [25:0] acqNet_io_out_2_bits_payload_addr_block;
  wire  acqNet_io_out_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_2_bits_payload_addr_beat;
  wire  acqNet_io_out_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_2_bits_payload_a_type;
  wire [10:0] acqNet_io_out_2_bits_payload_union;
  wire [63:0] acqNet_io_out_2_bits_payload_data;
  wire  acqNet_io_out_3_ready;
  wire  acqNet_io_out_3_valid;
  wire [1:0] acqNet_io_out_3_bits_header_src;
  wire [1:0] acqNet_io_out_3_bits_header_dst;
  wire [25:0] acqNet_io_out_3_bits_payload_addr_block;
  wire  acqNet_io_out_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_3_bits_payload_addr_beat;
  wire  acqNet_io_out_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_3_bits_payload_a_type;
  wire [10:0] acqNet_io_out_3_bits_payload_union;
  wire [63:0] acqNet_io_out_3_bits_payload_data;
  wire  relNet_clk;
  wire  relNet_reset;
  wire  relNet_io_in_0_ready;
  wire  relNet_io_in_0_valid;
  wire [1:0] relNet_io_in_0_bits_header_src;
  wire [1:0] relNet_io_in_0_bits_header_dst;
  wire [2:0] relNet_io_in_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_0_bits_payload_addr_block;
  wire  relNet_io_in_0_bits_payload_client_xact_id;
  wire  relNet_io_in_0_bits_payload_voluntary;
  wire [2:0] relNet_io_in_0_bits_payload_r_type;
  wire [63:0] relNet_io_in_0_bits_payload_data;
  wire  relNet_io_in_1_ready;
  wire  relNet_io_in_1_valid;
  wire [1:0] relNet_io_in_1_bits_header_src;
  wire [1:0] relNet_io_in_1_bits_header_dst;
  wire [2:0] relNet_io_in_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_1_bits_payload_addr_block;
  wire  relNet_io_in_1_bits_payload_client_xact_id;
  wire  relNet_io_in_1_bits_payload_voluntary;
  wire [2:0] relNet_io_in_1_bits_payload_r_type;
  wire [63:0] relNet_io_in_1_bits_payload_data;
  wire  relNet_io_in_2_ready;
  wire  relNet_io_in_2_valid;
  wire [1:0] relNet_io_in_2_bits_header_src;
  wire [1:0] relNet_io_in_2_bits_header_dst;
  wire [2:0] relNet_io_in_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_2_bits_payload_addr_block;
  wire  relNet_io_in_2_bits_payload_client_xact_id;
  wire  relNet_io_in_2_bits_payload_voluntary;
  wire [2:0] relNet_io_in_2_bits_payload_r_type;
  wire [63:0] relNet_io_in_2_bits_payload_data;
  wire  relNet_io_in_3_ready;
  wire  relNet_io_in_3_valid;
  wire [1:0] relNet_io_in_3_bits_header_src;
  wire [1:0] relNet_io_in_3_bits_header_dst;
  wire [2:0] relNet_io_in_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_3_bits_payload_addr_block;
  wire  relNet_io_in_3_bits_payload_client_xact_id;
  wire  relNet_io_in_3_bits_payload_voluntary;
  wire [2:0] relNet_io_in_3_bits_payload_r_type;
  wire [63:0] relNet_io_in_3_bits_payload_data;
  wire  relNet_io_out_0_ready;
  wire  relNet_io_out_0_valid;
  wire [1:0] relNet_io_out_0_bits_header_src;
  wire [1:0] relNet_io_out_0_bits_header_dst;
  wire [2:0] relNet_io_out_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_0_bits_payload_addr_block;
  wire  relNet_io_out_0_bits_payload_client_xact_id;
  wire  relNet_io_out_0_bits_payload_voluntary;
  wire [2:0] relNet_io_out_0_bits_payload_r_type;
  wire [63:0] relNet_io_out_0_bits_payload_data;
  wire  relNet_io_out_1_ready;
  wire  relNet_io_out_1_valid;
  wire [1:0] relNet_io_out_1_bits_header_src;
  wire [1:0] relNet_io_out_1_bits_header_dst;
  wire [2:0] relNet_io_out_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_1_bits_payload_addr_block;
  wire  relNet_io_out_1_bits_payload_client_xact_id;
  wire  relNet_io_out_1_bits_payload_voluntary;
  wire [2:0] relNet_io_out_1_bits_payload_r_type;
  wire [63:0] relNet_io_out_1_bits_payload_data;
  wire  relNet_io_out_2_ready;
  wire  relNet_io_out_2_valid;
  wire [1:0] relNet_io_out_2_bits_header_src;
  wire [1:0] relNet_io_out_2_bits_header_dst;
  wire [2:0] relNet_io_out_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_2_bits_payload_addr_block;
  wire  relNet_io_out_2_bits_payload_client_xact_id;
  wire  relNet_io_out_2_bits_payload_voluntary;
  wire [2:0] relNet_io_out_2_bits_payload_r_type;
  wire [63:0] relNet_io_out_2_bits_payload_data;
  wire  relNet_io_out_3_ready;
  wire  relNet_io_out_3_valid;
  wire [1:0] relNet_io_out_3_bits_header_src;
  wire [1:0] relNet_io_out_3_bits_header_dst;
  wire [2:0] relNet_io_out_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_3_bits_payload_addr_block;
  wire  relNet_io_out_3_bits_payload_client_xact_id;
  wire  relNet_io_out_3_bits_payload_voluntary;
  wire [2:0] relNet_io_out_3_bits_payload_r_type;
  wire [63:0] relNet_io_out_3_bits_payload_data;
  wire  prbNet_clk;
  wire  prbNet_reset;
  wire  prbNet_io_in_0_ready;
  wire  prbNet_io_in_0_valid;
  wire [1:0] prbNet_io_in_0_bits_header_src;
  wire [1:0] prbNet_io_in_0_bits_header_dst;
  wire [25:0] prbNet_io_in_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_0_bits_payload_p_type;
  wire  prbNet_io_in_1_ready;
  wire  prbNet_io_in_1_valid;
  wire [1:0] prbNet_io_in_1_bits_header_src;
  wire [1:0] prbNet_io_in_1_bits_header_dst;
  wire [25:0] prbNet_io_in_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_1_bits_payload_p_type;
  wire  prbNet_io_in_2_ready;
  wire  prbNet_io_in_2_valid;
  wire [1:0] prbNet_io_in_2_bits_header_src;
  wire [1:0] prbNet_io_in_2_bits_header_dst;
  wire [25:0] prbNet_io_in_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_2_bits_payload_p_type;
  wire  prbNet_io_in_3_ready;
  wire  prbNet_io_in_3_valid;
  wire [1:0] prbNet_io_in_3_bits_header_src;
  wire [1:0] prbNet_io_in_3_bits_header_dst;
  wire [25:0] prbNet_io_in_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_3_bits_payload_p_type;
  wire  prbNet_io_out_0_ready;
  wire  prbNet_io_out_0_valid;
  wire [1:0] prbNet_io_out_0_bits_header_src;
  wire [1:0] prbNet_io_out_0_bits_header_dst;
  wire [25:0] prbNet_io_out_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_0_bits_payload_p_type;
  wire  prbNet_io_out_1_ready;
  wire  prbNet_io_out_1_valid;
  wire [1:0] prbNet_io_out_1_bits_header_src;
  wire [1:0] prbNet_io_out_1_bits_header_dst;
  wire [25:0] prbNet_io_out_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_1_bits_payload_p_type;
  wire  prbNet_io_out_2_ready;
  wire  prbNet_io_out_2_valid;
  wire [1:0] prbNet_io_out_2_bits_header_src;
  wire [1:0] prbNet_io_out_2_bits_header_dst;
  wire [25:0] prbNet_io_out_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_2_bits_payload_p_type;
  wire  prbNet_io_out_3_ready;
  wire  prbNet_io_out_3_valid;
  wire [1:0] prbNet_io_out_3_bits_header_src;
  wire [1:0] prbNet_io_out_3_bits_header_dst;
  wire [25:0] prbNet_io_out_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_3_bits_payload_p_type;
  wire  gntNet_clk;
  wire  gntNet_reset;
  wire  gntNet_io_in_0_ready;
  wire  gntNet_io_in_0_valid;
  wire [1:0] gntNet_io_in_0_bits_header_src;
  wire [1:0] gntNet_io_in_0_bits_header_dst;
  wire [2:0] gntNet_io_in_0_bits_payload_addr_beat;
  wire  gntNet_io_in_0_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_in_0_bits_payload_manager_xact_id;
  wire  gntNet_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_0_bits_payload_g_type;
  wire [63:0] gntNet_io_in_0_bits_payload_data;
  wire  gntNet_io_in_1_ready;
  wire  gntNet_io_in_1_valid;
  wire [1:0] gntNet_io_in_1_bits_header_src;
  wire [1:0] gntNet_io_in_1_bits_header_dst;
  wire [2:0] gntNet_io_in_1_bits_payload_addr_beat;
  wire  gntNet_io_in_1_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_in_1_bits_payload_manager_xact_id;
  wire  gntNet_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_1_bits_payload_g_type;
  wire [63:0] gntNet_io_in_1_bits_payload_data;
  wire  gntNet_io_in_2_ready;
  wire  gntNet_io_in_2_valid;
  wire [1:0] gntNet_io_in_2_bits_header_src;
  wire [1:0] gntNet_io_in_2_bits_header_dst;
  wire [2:0] gntNet_io_in_2_bits_payload_addr_beat;
  wire  gntNet_io_in_2_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_in_2_bits_payload_manager_xact_id;
  wire  gntNet_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_2_bits_payload_g_type;
  wire [63:0] gntNet_io_in_2_bits_payload_data;
  wire  gntNet_io_in_3_ready;
  wire  gntNet_io_in_3_valid;
  wire [1:0] gntNet_io_in_3_bits_header_src;
  wire [1:0] gntNet_io_in_3_bits_header_dst;
  wire [2:0] gntNet_io_in_3_bits_payload_addr_beat;
  wire  gntNet_io_in_3_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_in_3_bits_payload_manager_xact_id;
  wire  gntNet_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_3_bits_payload_g_type;
  wire [63:0] gntNet_io_in_3_bits_payload_data;
  wire  gntNet_io_out_0_ready;
  wire  gntNet_io_out_0_valid;
  wire [1:0] gntNet_io_out_0_bits_header_src;
  wire [1:0] gntNet_io_out_0_bits_header_dst;
  wire [2:0] gntNet_io_out_0_bits_payload_addr_beat;
  wire  gntNet_io_out_0_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_out_0_bits_payload_manager_xact_id;
  wire  gntNet_io_out_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_0_bits_payload_g_type;
  wire [63:0] gntNet_io_out_0_bits_payload_data;
  wire  gntNet_io_out_1_ready;
  wire  gntNet_io_out_1_valid;
  wire [1:0] gntNet_io_out_1_bits_header_src;
  wire [1:0] gntNet_io_out_1_bits_header_dst;
  wire [2:0] gntNet_io_out_1_bits_payload_addr_beat;
  wire  gntNet_io_out_1_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_out_1_bits_payload_manager_xact_id;
  wire  gntNet_io_out_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_1_bits_payload_g_type;
  wire [63:0] gntNet_io_out_1_bits_payload_data;
  wire  gntNet_io_out_2_ready;
  wire  gntNet_io_out_2_valid;
  wire [1:0] gntNet_io_out_2_bits_header_src;
  wire [1:0] gntNet_io_out_2_bits_header_dst;
  wire [2:0] gntNet_io_out_2_bits_payload_addr_beat;
  wire  gntNet_io_out_2_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_out_2_bits_payload_manager_xact_id;
  wire  gntNet_io_out_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_2_bits_payload_g_type;
  wire [63:0] gntNet_io_out_2_bits_payload_data;
  wire  gntNet_io_out_3_ready;
  wire  gntNet_io_out_3_valid;
  wire [1:0] gntNet_io_out_3_bits_header_src;
  wire [1:0] gntNet_io_out_3_bits_header_dst;
  wire [2:0] gntNet_io_out_3_bits_payload_addr_beat;
  wire  gntNet_io_out_3_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_out_3_bits_payload_manager_xact_id;
  wire  gntNet_io_out_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_3_bits_payload_g_type;
  wire [63:0] gntNet_io_out_3_bits_payload_data;
  wire  ackNet_clk;
  wire  ackNet_reset;
  wire  ackNet_io_in_0_ready;
  wire  ackNet_io_in_0_valid;
  wire [1:0] ackNet_io_in_0_bits_header_src;
  wire [1:0] ackNet_io_in_0_bits_header_dst;
  wire [1:0] ackNet_io_in_0_bits_payload_manager_xact_id;
  wire  ackNet_io_in_1_ready;
  wire  ackNet_io_in_1_valid;
  wire [1:0] ackNet_io_in_1_bits_header_src;
  wire [1:0] ackNet_io_in_1_bits_header_dst;
  wire [1:0] ackNet_io_in_1_bits_payload_manager_xact_id;
  wire  ackNet_io_in_2_ready;
  wire  ackNet_io_in_2_valid;
  wire [1:0] ackNet_io_in_2_bits_header_src;
  wire [1:0] ackNet_io_in_2_bits_header_dst;
  wire [1:0] ackNet_io_in_2_bits_payload_manager_xact_id;
  wire  ackNet_io_in_3_ready;
  wire  ackNet_io_in_3_valid;
  wire [1:0] ackNet_io_in_3_bits_header_src;
  wire [1:0] ackNet_io_in_3_bits_header_dst;
  wire [1:0] ackNet_io_in_3_bits_payload_manager_xact_id;
  wire  ackNet_io_out_0_ready;
  wire  ackNet_io_out_0_valid;
  wire [1:0] ackNet_io_out_0_bits_header_src;
  wire [1:0] ackNet_io_out_0_bits_header_dst;
  wire [1:0] ackNet_io_out_0_bits_payload_manager_xact_id;
  wire  ackNet_io_out_1_ready;
  wire  ackNet_io_out_1_valid;
  wire [1:0] ackNet_io_out_1_bits_header_src;
  wire [1:0] ackNet_io_out_1_bits_header_dst;
  wire [1:0] ackNet_io_out_1_bits_payload_manager_xact_id;
  wire  ackNet_io_out_2_ready;
  wire  ackNet_io_out_2_valid;
  wire [1:0] ackNet_io_out_2_bits_header_src;
  wire [1:0] ackNet_io_out_2_bits_header_dst;
  wire [1:0] ackNet_io_out_2_bits_payload_manager_xact_id;
  wire  ackNet_io_out_3_ready;
  wire  ackNet_io_out_3_valid;
  wire [1:0] ackNet_io_out_3_bits_header_src;
  wire [1:0] ackNet_io_out_3_bits_header_dst;
  wire [1:0] ackNet_io_out_3_bits_payload_manager_xact_id;
  wire  T_12724_ready;
  wire  T_12724_valid;
  wire [1:0] T_12724_bits_header_src;
  wire [1:0] T_12724_bits_header_dst;
  wire [25:0] T_12724_bits_payload_addr_block;
  wire  T_12724_bits_payload_client_xact_id;
  wire [2:0] T_12724_bits_payload_addr_beat;
  wire  T_12724_bits_payload_is_builtin_type;
  wire [2:0] T_12724_bits_payload_a_type;
  wire [10:0] T_12724_bits_payload_union;
  wire [63:0] T_12724_bits_payload_data;
  wire [2:0] T_12952;
  wire [1:0] T_12953;
  wire  T_13294_ready;
  wire  T_13294_valid;
  wire [1:0] T_13294_bits_header_src;
  wire [1:0] T_13294_bits_header_dst;
  wire [25:0] T_13294_bits_payload_addr_block;
  wire  T_13294_bits_payload_client_xact_id;
  wire [2:0] T_13294_bits_payload_addr_beat;
  wire  T_13294_bits_payload_is_builtin_type;
  wire [2:0] T_13294_bits_payload_a_type;
  wire [10:0] T_13294_bits_payload_union;
  wire [63:0] T_13294_bits_payload_data;
  wire [2:0] T_13522;
  wire [1:0] T_13523;
  wire  T_13624_ready;
  wire  T_13624_valid;
  wire [1:0] T_13624_bits_header_src;
  wire [1:0] T_13624_bits_header_dst;
  wire [25:0] T_13624_bits_payload_addr_block;
  wire  T_13624_bits_payload_client_xact_id;
  wire [2:0] T_13624_bits_payload_addr_beat;
  wire  T_13624_bits_payload_is_builtin_type;
  wire [2:0] T_13624_bits_payload_a_type;
  wire [10:0] T_13624_bits_payload_union;
  wire [63:0] T_13624_bits_payload_data;
  wire [2:0] T_13692;
  wire [1:0] T_13693;
  wire  T_13794_ready;
  wire  T_13794_valid;
  wire [1:0] T_13794_bits_header_src;
  wire [1:0] T_13794_bits_header_dst;
  wire [25:0] T_13794_bits_payload_addr_block;
  wire  T_13794_bits_payload_client_xact_id;
  wire [2:0] T_13794_bits_payload_addr_beat;
  wire  T_13794_bits_payload_is_builtin_type;
  wire [2:0] T_13794_bits_payload_a_type;
  wire [10:0] T_13794_bits_payload_union;
  wire [63:0] T_13794_bits_payload_data;
  wire [2:0] T_13862;
  wire [1:0] T_13863;
  wire  T_14201_ready;
  wire  T_14201_valid;
  wire [1:0] T_14201_bits_header_src;
  wire [1:0] T_14201_bits_header_dst;
  wire [2:0] T_14201_bits_payload_addr_beat;
  wire [25:0] T_14201_bits_payload_addr_block;
  wire  T_14201_bits_payload_client_xact_id;
  wire  T_14201_bits_payload_voluntary;
  wire [2:0] T_14201_bits_payload_r_type;
  wire [63:0] T_14201_bits_payload_data;
  wire [2:0] T_14427;
  wire [1:0] T_14428;
  wire  T_14766_ready;
  wire  T_14766_valid;
  wire [1:0] T_14766_bits_header_src;
  wire [1:0] T_14766_bits_header_dst;
  wire [2:0] T_14766_bits_payload_addr_beat;
  wire [25:0] T_14766_bits_payload_addr_block;
  wire  T_14766_bits_payload_client_xact_id;
  wire  T_14766_bits_payload_voluntary;
  wire [2:0] T_14766_bits_payload_r_type;
  wire [63:0] T_14766_bits_payload_data;
  wire [2:0] T_14992;
  wire [1:0] T_14993;
  wire  T_15091_ready;
  wire  T_15091_valid;
  wire [1:0] T_15091_bits_header_src;
  wire [1:0] T_15091_bits_header_dst;
  wire [2:0] T_15091_bits_payload_addr_beat;
  wire [25:0] T_15091_bits_payload_addr_block;
  wire  T_15091_bits_payload_client_xact_id;
  wire  T_15091_bits_payload_voluntary;
  wire [2:0] T_15091_bits_payload_r_type;
  wire [63:0] T_15091_bits_payload_data;
  wire [2:0] T_15157;
  wire [1:0] T_15158;
  wire  T_15256_ready;
  wire  T_15256_valid;
  wire [1:0] T_15256_bits_header_src;
  wire [1:0] T_15256_bits_header_dst;
  wire [2:0] T_15256_bits_payload_addr_beat;
  wire [25:0] T_15256_bits_payload_addr_block;
  wire  T_15256_bits_payload_client_xact_id;
  wire  T_15256_bits_payload_voluntary;
  wire [2:0] T_15256_bits_payload_r_type;
  wire [63:0] T_15256_bits_payload_data;
  wire [2:0] T_15322;
  wire [1:0] T_15323;
  wire  T_15409_ready;
  wire  T_15409_valid;
  wire [1:0] T_15409_bits_header_src;
  wire [1:0] T_15409_bits_header_dst;
  wire [25:0] T_15409_bits_payload_addr_block;
  wire [1:0] T_15409_bits_payload_p_type;
  wire [2:0] T_15467;
  wire [1:0] T_15468;
  wire  T_15554_ready;
  wire  T_15554_valid;
  wire [1:0] T_15554_bits_header_src;
  wire [1:0] T_15554_bits_header_dst;
  wire [25:0] T_15554_bits_payload_addr_block;
  wire [1:0] T_15554_bits_payload_p_type;
  wire [2:0] T_15612;
  wire [1:0] T_15613;
  wire  T_15939_ready;
  wire  T_15939_valid;
  wire [1:0] T_15939_bits_header_src;
  wire [1:0] T_15939_bits_header_dst;
  wire [25:0] T_15939_bits_payload_addr_block;
  wire [1:0] T_15939_bits_payload_p_type;
  wire [2:0] T_16157;
  wire [1:0] T_16158;
  wire  T_16484_ready;
  wire  T_16484_valid;
  wire [1:0] T_16484_bits_header_src;
  wire [1:0] T_16484_bits_header_dst;
  wire [25:0] T_16484_bits_payload_addr_block;
  wire [1:0] T_16484_bits_payload_p_type;
  wire [2:0] T_16702;
  wire [1:0] T_16703;
  wire  T_16801_ready;
  wire  T_16801_valid;
  wire [1:0] T_16801_bits_header_src;
  wire [1:0] T_16801_bits_header_dst;
  wire [2:0] T_16801_bits_payload_addr_beat;
  wire  T_16801_bits_payload_client_xact_id;
  wire [1:0] T_16801_bits_payload_manager_xact_id;
  wire  T_16801_bits_payload_is_builtin_type;
  wire [3:0] T_16801_bits_payload_g_type;
  wire [63:0] T_16801_bits_payload_data;
  wire [2:0] T_16867;
  wire [1:0] T_16868;
  wire  T_16966_ready;
  wire  T_16966_valid;
  wire [1:0] T_16966_bits_header_src;
  wire [1:0] T_16966_bits_header_dst;
  wire [2:0] T_16966_bits_payload_addr_beat;
  wire  T_16966_bits_payload_client_xact_id;
  wire [1:0] T_16966_bits_payload_manager_xact_id;
  wire  T_16966_bits_payload_is_builtin_type;
  wire [3:0] T_16966_bits_payload_g_type;
  wire [63:0] T_16966_bits_payload_data;
  wire [2:0] T_17032;
  wire [1:0] T_17033;
  wire  T_17371_ready;
  wire  T_17371_valid;
  wire [1:0] T_17371_bits_header_src;
  wire [1:0] T_17371_bits_header_dst;
  wire [2:0] T_17371_bits_payload_addr_beat;
  wire  T_17371_bits_payload_client_xact_id;
  wire [1:0] T_17371_bits_payload_manager_xact_id;
  wire  T_17371_bits_payload_is_builtin_type;
  wire [3:0] T_17371_bits_payload_g_type;
  wire [63:0] T_17371_bits_payload_data;
  wire [2:0] T_17597;
  wire [1:0] T_17598;
  wire  T_17936_ready;
  wire  T_17936_valid;
  wire [1:0] T_17936_bits_header_src;
  wire [1:0] T_17936_bits_header_dst;
  wire [2:0] T_17936_bits_payload_addr_beat;
  wire  T_17936_bits_payload_client_xact_id;
  wire [1:0] T_17936_bits_payload_manager_xact_id;
  wire  T_17936_bits_payload_is_builtin_type;
  wire [3:0] T_17936_bits_payload_g_type;
  wire [63:0] T_17936_bits_payload_data;
  wire [2:0] T_18162;
  wire [1:0] T_18163;
  wire  T_18486_ready;
  wire  T_18486_valid;
  wire [1:0] T_18486_bits_header_src;
  wire [1:0] T_18486_bits_header_dst;
  wire [1:0] T_18486_bits_payload_manager_xact_id;
  wire [2:0] T_18702;
  wire [1:0] T_18703;
  wire  T_19026_ready;
  wire  T_19026_valid;
  wire [1:0] T_19026_bits_header_src;
  wire [1:0] T_19026_bits_header_dst;
  wire [1:0] T_19026_bits_payload_manager_xact_id;
  wire [2:0] T_19242;
  wire [1:0] T_19243;
  wire  T_19326_ready;
  wire  T_19326_valid;
  wire [1:0] T_19326_bits_header_src;
  wire [1:0] T_19326_bits_header_dst;
  wire [1:0] T_19326_bits_payload_manager_xact_id;
  wire [2:0] T_19382;
  wire [1:0] T_19383;
  wire  T_19466_ready;
  wire  T_19466_valid;
  wire [1:0] T_19466_bits_header_src;
  wire [1:0] T_19466_bits_header_dst;
  wire [1:0] T_19466_bits_payload_manager_xact_id;
  wire [2:0] T_19522;
  wire [1:0] T_19523;
  wire [1:0] GEN_0;
  reg [31:0] GEN_64;
  wire [1:0] GEN_1;
  reg [31:0] GEN_65;
  wire [25:0] GEN_2;
  reg [31:0] GEN_66;
  wire  GEN_3;
  reg [31:0] GEN_67;
  wire [2:0] GEN_4;
  reg [31:0] GEN_68;
  wire  GEN_5;
  reg [31:0] GEN_69;
  wire [2:0] GEN_6;
  reg [31:0] GEN_70;
  wire [10:0] GEN_7;
  reg [31:0] GEN_71;
  wire [63:0] GEN_8;
  reg [63:0] GEN_72;
  wire [1:0] GEN_9;
  reg [31:0] GEN_73;
  wire [1:0] GEN_10;
  reg [31:0] GEN_74;
  wire [25:0] GEN_11;
  reg [31:0] GEN_75;
  wire  GEN_12;
  reg [31:0] GEN_76;
  wire [2:0] GEN_13;
  reg [31:0] GEN_77;
  wire  GEN_14;
  reg [31:0] GEN_78;
  wire [2:0] GEN_15;
  reg [31:0] GEN_79;
  wire [10:0] GEN_16;
  reg [31:0] GEN_80;
  wire [63:0] GEN_17;
  reg [63:0] GEN_81;
  wire [1:0] GEN_18;
  reg [31:0] GEN_82;
  wire [1:0] GEN_19;
  reg [31:0] GEN_83;
  wire [2:0] GEN_20;
  reg [31:0] GEN_84;
  wire [25:0] GEN_21;
  reg [31:0] GEN_85;
  wire  GEN_22;
  reg [31:0] GEN_86;
  wire  GEN_23;
  reg [31:0] GEN_87;
  wire [2:0] GEN_24;
  reg [31:0] GEN_88;
  wire [63:0] GEN_25;
  reg [63:0] GEN_89;
  wire [1:0] GEN_26;
  reg [31:0] GEN_90;
  wire [1:0] GEN_27;
  reg [31:0] GEN_91;
  wire [2:0] GEN_28;
  reg [31:0] GEN_92;
  wire [25:0] GEN_29;
  reg [31:0] GEN_93;
  wire  GEN_30;
  reg [31:0] GEN_94;
  wire  GEN_31;
  reg [31:0] GEN_95;
  wire [2:0] GEN_32;
  reg [31:0] GEN_96;
  wire [63:0] GEN_33;
  reg [63:0] GEN_97;
  wire [1:0] GEN_34;
  reg [31:0] GEN_98;
  wire [1:0] GEN_35;
  reg [31:0] GEN_99;
  wire [25:0] GEN_36;
  reg [31:0] GEN_100;
  wire [1:0] GEN_37;
  reg [31:0] GEN_101;
  wire [1:0] GEN_38;
  reg [31:0] GEN_102;
  wire [1:0] GEN_39;
  reg [31:0] GEN_103;
  wire [25:0] GEN_40;
  reg [31:0] GEN_104;
  wire [1:0] GEN_41;
  reg [31:0] GEN_105;
  wire [1:0] GEN_42;
  reg [31:0] GEN_106;
  wire [1:0] GEN_43;
  reg [31:0] GEN_107;
  wire [2:0] GEN_44;
  reg [31:0] GEN_108;
  wire  GEN_45;
  reg [31:0] GEN_109;
  wire [1:0] GEN_46;
  reg [31:0] GEN_110;
  wire  GEN_47;
  reg [31:0] GEN_111;
  wire [3:0] GEN_48;
  reg [31:0] GEN_112;
  wire [63:0] GEN_49;
  reg [63:0] GEN_113;
  wire [1:0] GEN_50;
  reg [31:0] GEN_114;
  wire [1:0] GEN_51;
  reg [31:0] GEN_115;
  wire [2:0] GEN_52;
  reg [31:0] GEN_116;
  wire  GEN_53;
  reg [31:0] GEN_117;
  wire [1:0] GEN_54;
  reg [31:0] GEN_118;
  wire  GEN_55;
  reg [31:0] GEN_119;
  wire [3:0] GEN_56;
  reg [31:0] GEN_120;
  wire [63:0] GEN_57;
  reg [63:0] GEN_121;
  wire [1:0] GEN_58;
  reg [31:0] GEN_122;
  wire [1:0] GEN_59;
  reg [31:0] GEN_123;
  wire [1:0] GEN_60;
  reg [31:0] GEN_124;
  wire [1:0] GEN_61;
  reg [31:0] GEN_125;
  wire [1:0] GEN_62;
  reg [31:0] GEN_126;
  wire [1:0] GEN_63;
  reg [31:0] GEN_127;
  TileLinkEnqueuer TileLinkEnqueuer_4 (
    .clk(TileLinkEnqueuer_4_clk),
    .reset(TileLinkEnqueuer_4_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_4_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_4_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_4_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_4_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_4_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_4_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_4_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_4_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_4_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_4_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_4_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_4_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_4_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_4_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_4_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_4_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_4_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_4_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_4_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_4_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_4_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_4_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_4_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_4_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_4_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_4_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_4_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_4_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_4_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_4_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_4_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_4_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_4_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_4_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_4_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_4_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_4_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_4_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_4_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_4_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_4_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_4_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_4_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_4_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_4_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_4_io_manager_release_bits_payload_data)
  );
  ClientTileLinkNetworkPort ClientTileLinkNetworkPort_1 (
    .clk(ClientTileLinkNetworkPort_1_clk),
    .reset(ClientTileLinkNetworkPort_1_reset),
    .io_client_acquire_ready(ClientTileLinkNetworkPort_1_io_client_acquire_ready),
    .io_client_acquire_valid(ClientTileLinkNetworkPort_1_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientTileLinkNetworkPort_1_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientTileLinkNetworkPort_1_io_client_acquire_bits_data),
    .io_client_probe_ready(ClientTileLinkNetworkPort_1_io_client_probe_ready),
    .io_client_probe_valid(ClientTileLinkNetworkPort_1_io_client_probe_valid),
    .io_client_probe_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block),
    .io_client_probe_bits_p_type(ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type),
    .io_client_release_ready(ClientTileLinkNetworkPort_1_io_client_release_ready),
    .io_client_release_valid(ClientTileLinkNetworkPort_1_io_client_release_valid),
    .io_client_release_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat),
    .io_client_release_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block),
    .io_client_release_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id),
    .io_client_release_bits_voluntary(ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary),
    .io_client_release_bits_r_type(ClientTileLinkNetworkPort_1_io_client_release_bits_r_type),
    .io_client_release_bits_data(ClientTileLinkNetworkPort_1_io_client_release_bits_data),
    .io_client_grant_ready(ClientTileLinkNetworkPort_1_io_client_grant_ready),
    .io_client_grant_valid(ClientTileLinkNetworkPort_1_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientTileLinkNetworkPort_1_io_client_grant_bits_data),
    .io_client_grant_bits_manager_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id),
    .io_client_finish_ready(ClientTileLinkNetworkPort_1_io_client_finish_ready),
    .io_client_finish_valid(ClientTileLinkNetworkPort_1_io_client_finish_valid),
    .io_client_finish_bits_manager_xact_id(ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id),
    .io_client_finish_bits_manager_id(ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id),
    .io_network_acquire_ready(ClientTileLinkNetworkPort_1_io_network_acquire_ready),
    .io_network_acquire_valid(ClientTileLinkNetworkPort_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientTileLinkNetworkPort_1_io_network_grant_ready),
    .io_network_grant_valid(ClientTileLinkNetworkPort_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientTileLinkNetworkPort_1_io_network_finish_ready),
    .io_network_finish_valid(ClientTileLinkNetworkPort_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientTileLinkNetworkPort_1_io_network_probe_ready),
    .io_network_probe_valid(ClientTileLinkNetworkPort_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientTileLinkNetworkPort_1_io_network_release_ready),
    .io_network_release_valid(ClientTileLinkNetworkPort_1_io_network_release_valid),
    .io_network_release_bits_header_src(ClientTileLinkNetworkPort_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_1_1 (
    .clk(TileLinkEnqueuer_1_1_clk),
    .reset(TileLinkEnqueuer_1_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_1_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_1_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_1_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_1_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_1_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_1_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_1_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_1_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_1_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_1_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_1_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_1_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_1_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_1_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_1_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_1_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_1_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_1_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_1_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_1_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_1_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_1_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_1_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_1_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_1_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_1_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_1_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data)
  );
  ClientUncachedTileLinkNetworkPort ClientUncachedTileLinkNetworkPort_1 (
    .clk(ClientUncachedTileLinkNetworkPort_1_clk),
    .reset(ClientUncachedTileLinkNetworkPort_1_reset),
    .io_client_acquire_ready(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready),
    .io_client_acquire_valid(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data),
    .io_client_grant_ready(ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready),
    .io_client_grant_valid(ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data),
    .io_network_acquire_ready(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready),
    .io_network_acquire_valid(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready),
    .io_network_grant_valid(ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready),
    .io_network_finish_valid(ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready),
    .io_network_probe_valid(ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientUncachedTileLinkNetworkPort_1_io_network_release_ready),
    .io_network_release_valid(ClientUncachedTileLinkNetworkPort_1_io_network_release_valid),
    .io_network_release_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort ManagerTileLinkNetworkPort_2 (
    .clk(ManagerTileLinkNetworkPort_2_clk),
    .reset(ManagerTileLinkNetworkPort_2_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_2_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_2_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_2_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_2_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_2_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_2_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_2_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_2_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_2_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_2_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_2_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_2_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_2_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_2_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_2_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_2_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_2_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_2_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_2_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_2_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_2_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_2 TileLinkEnqueuer_2_1 (
    .clk(TileLinkEnqueuer_2_1_clk),
    .reset(TileLinkEnqueuer_2_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_2_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_2_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_2_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_2_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_2_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_2_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_2_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_2_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_2_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_2_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_2_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_2_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_2_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_2_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_2_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_2_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_2_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_2_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_2_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_2_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_2_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_2_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_2_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_2_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_2_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_2_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_2_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort_1 ManagerTileLinkNetworkPort_1_1 (
    .clk(ManagerTileLinkNetworkPort_1_1_clk),
    .reset(ManagerTileLinkNetworkPort_1_1_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_1_1_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_1_1_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_1_1_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_1_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_1_1_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_1_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_1_1_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_1_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_1_1_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_1_1_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_2 TileLinkEnqueuer_3_1 (
    .clk(TileLinkEnqueuer_3_1_clk),
    .reset(TileLinkEnqueuer_3_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_3_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_3_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_3_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_3_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_3_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_3_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_3_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_3_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_3_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_3_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_3_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_3_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_3_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_3_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_3_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_3_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_3_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_3_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_3_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_3_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_3_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_3_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_3_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_3_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_3_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_3_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_3_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data)
  );
  BasicBus acqNet (
    .clk(acqNet_clk),
    .reset(acqNet_reset),
    .io_in_0_ready(acqNet_io_in_0_ready),
    .io_in_0_valid(acqNet_io_in_0_valid),
    .io_in_0_bits_header_src(acqNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(acqNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(acqNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(acqNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(acqNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(acqNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(acqNet_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(acqNet_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(acqNet_io_in_0_bits_payload_data),
    .io_in_1_ready(acqNet_io_in_1_ready),
    .io_in_1_valid(acqNet_io_in_1_valid),
    .io_in_1_bits_header_src(acqNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(acqNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(acqNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(acqNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(acqNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(acqNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(acqNet_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(acqNet_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(acqNet_io_in_1_bits_payload_data),
    .io_in_2_ready(acqNet_io_in_2_ready),
    .io_in_2_valid(acqNet_io_in_2_valid),
    .io_in_2_bits_header_src(acqNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(acqNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(acqNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(acqNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(acqNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(acqNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(acqNet_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(acqNet_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(acqNet_io_in_2_bits_payload_data),
    .io_in_3_ready(acqNet_io_in_3_ready),
    .io_in_3_valid(acqNet_io_in_3_valid),
    .io_in_3_bits_header_src(acqNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(acqNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(acqNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(acqNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(acqNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(acqNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(acqNet_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(acqNet_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(acqNet_io_in_3_bits_payload_data),
    .io_out_0_ready(acqNet_io_out_0_ready),
    .io_out_0_valid(acqNet_io_out_0_valid),
    .io_out_0_bits_header_src(acqNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(acqNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(acqNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(acqNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_addr_beat(acqNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_is_builtin_type(acqNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_a_type(acqNet_io_out_0_bits_payload_a_type),
    .io_out_0_bits_payload_union(acqNet_io_out_0_bits_payload_union),
    .io_out_0_bits_payload_data(acqNet_io_out_0_bits_payload_data),
    .io_out_1_ready(acqNet_io_out_1_ready),
    .io_out_1_valid(acqNet_io_out_1_valid),
    .io_out_1_bits_header_src(acqNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(acqNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(acqNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(acqNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_addr_beat(acqNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_is_builtin_type(acqNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_a_type(acqNet_io_out_1_bits_payload_a_type),
    .io_out_1_bits_payload_union(acqNet_io_out_1_bits_payload_union),
    .io_out_1_bits_payload_data(acqNet_io_out_1_bits_payload_data),
    .io_out_2_ready(acqNet_io_out_2_ready),
    .io_out_2_valid(acqNet_io_out_2_valid),
    .io_out_2_bits_header_src(acqNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(acqNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(acqNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(acqNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_addr_beat(acqNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_is_builtin_type(acqNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_a_type(acqNet_io_out_2_bits_payload_a_type),
    .io_out_2_bits_payload_union(acqNet_io_out_2_bits_payload_union),
    .io_out_2_bits_payload_data(acqNet_io_out_2_bits_payload_data),
    .io_out_3_ready(acqNet_io_out_3_ready),
    .io_out_3_valid(acqNet_io_out_3_valid),
    .io_out_3_bits_header_src(acqNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(acqNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(acqNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(acqNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_addr_beat(acqNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_is_builtin_type(acqNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_a_type(acqNet_io_out_3_bits_payload_a_type),
    .io_out_3_bits_payload_union(acqNet_io_out_3_bits_payload_union),
    .io_out_3_bits_payload_data(acqNet_io_out_3_bits_payload_data)
  );
  BasicBus_1 relNet (
    .clk(relNet_clk),
    .reset(relNet_reset),
    .io_in_0_ready(relNet_io_in_0_ready),
    .io_in_0_valid(relNet_io_in_0_valid),
    .io_in_0_bits_header_src(relNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(relNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(relNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(relNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(relNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(relNet_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(relNet_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(relNet_io_in_0_bits_payload_data),
    .io_in_1_ready(relNet_io_in_1_ready),
    .io_in_1_valid(relNet_io_in_1_valid),
    .io_in_1_bits_header_src(relNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(relNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(relNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(relNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(relNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(relNet_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(relNet_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(relNet_io_in_1_bits_payload_data),
    .io_in_2_ready(relNet_io_in_2_ready),
    .io_in_2_valid(relNet_io_in_2_valid),
    .io_in_2_bits_header_src(relNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(relNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(relNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(relNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(relNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(relNet_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(relNet_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(relNet_io_in_2_bits_payload_data),
    .io_in_3_ready(relNet_io_in_3_ready),
    .io_in_3_valid(relNet_io_in_3_valid),
    .io_in_3_bits_header_src(relNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(relNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(relNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(relNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(relNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(relNet_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(relNet_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(relNet_io_in_3_bits_payload_data),
    .io_out_0_ready(relNet_io_out_0_ready),
    .io_out_0_valid(relNet_io_out_0_valid),
    .io_out_0_bits_header_src(relNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(relNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(relNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_addr_block(relNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(relNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_voluntary(relNet_io_out_0_bits_payload_voluntary),
    .io_out_0_bits_payload_r_type(relNet_io_out_0_bits_payload_r_type),
    .io_out_0_bits_payload_data(relNet_io_out_0_bits_payload_data),
    .io_out_1_ready(relNet_io_out_1_ready),
    .io_out_1_valid(relNet_io_out_1_valid),
    .io_out_1_bits_header_src(relNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(relNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(relNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_addr_block(relNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(relNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_voluntary(relNet_io_out_1_bits_payload_voluntary),
    .io_out_1_bits_payload_r_type(relNet_io_out_1_bits_payload_r_type),
    .io_out_1_bits_payload_data(relNet_io_out_1_bits_payload_data),
    .io_out_2_ready(relNet_io_out_2_ready),
    .io_out_2_valid(relNet_io_out_2_valid),
    .io_out_2_bits_header_src(relNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(relNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(relNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_addr_block(relNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(relNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_voluntary(relNet_io_out_2_bits_payload_voluntary),
    .io_out_2_bits_payload_r_type(relNet_io_out_2_bits_payload_r_type),
    .io_out_2_bits_payload_data(relNet_io_out_2_bits_payload_data),
    .io_out_3_ready(relNet_io_out_3_ready),
    .io_out_3_valid(relNet_io_out_3_valid),
    .io_out_3_bits_header_src(relNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(relNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(relNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_addr_block(relNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(relNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_voluntary(relNet_io_out_3_bits_payload_voluntary),
    .io_out_3_bits_payload_r_type(relNet_io_out_3_bits_payload_r_type),
    .io_out_3_bits_payload_data(relNet_io_out_3_bits_payload_data)
  );
  BasicBus_2 prbNet (
    .clk(prbNet_clk),
    .reset(prbNet_reset),
    .io_in_0_ready(prbNet_io_in_0_ready),
    .io_in_0_valid(prbNet_io_in_0_valid),
    .io_in_0_bits_header_src(prbNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(prbNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(prbNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(prbNet_io_in_0_bits_payload_p_type),
    .io_in_1_ready(prbNet_io_in_1_ready),
    .io_in_1_valid(prbNet_io_in_1_valid),
    .io_in_1_bits_header_src(prbNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(prbNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(prbNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(prbNet_io_in_1_bits_payload_p_type),
    .io_in_2_ready(prbNet_io_in_2_ready),
    .io_in_2_valid(prbNet_io_in_2_valid),
    .io_in_2_bits_header_src(prbNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(prbNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(prbNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(prbNet_io_in_2_bits_payload_p_type),
    .io_in_3_ready(prbNet_io_in_3_ready),
    .io_in_3_valid(prbNet_io_in_3_valid),
    .io_in_3_bits_header_src(prbNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(prbNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(prbNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(prbNet_io_in_3_bits_payload_p_type),
    .io_out_0_ready(prbNet_io_out_0_ready),
    .io_out_0_valid(prbNet_io_out_0_valid),
    .io_out_0_bits_header_src(prbNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(prbNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(prbNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_p_type(prbNet_io_out_0_bits_payload_p_type),
    .io_out_1_ready(prbNet_io_out_1_ready),
    .io_out_1_valid(prbNet_io_out_1_valid),
    .io_out_1_bits_header_src(prbNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(prbNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(prbNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_p_type(prbNet_io_out_1_bits_payload_p_type),
    .io_out_2_ready(prbNet_io_out_2_ready),
    .io_out_2_valid(prbNet_io_out_2_valid),
    .io_out_2_bits_header_src(prbNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(prbNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(prbNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_p_type(prbNet_io_out_2_bits_payload_p_type),
    .io_out_3_ready(prbNet_io_out_3_ready),
    .io_out_3_valid(prbNet_io_out_3_valid),
    .io_out_3_bits_header_src(prbNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(prbNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(prbNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_p_type(prbNet_io_out_3_bits_payload_p_type)
  );
  BasicBus_3 gntNet (
    .clk(gntNet_clk),
    .reset(gntNet_reset),
    .io_in_0_ready(gntNet_io_in_0_ready),
    .io_in_0_valid(gntNet_io_in_0_valid),
    .io_in_0_bits_header_src(gntNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(gntNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(gntNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(gntNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(gntNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(gntNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(gntNet_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(gntNet_io_in_0_bits_payload_data),
    .io_in_1_ready(gntNet_io_in_1_ready),
    .io_in_1_valid(gntNet_io_in_1_valid),
    .io_in_1_bits_header_src(gntNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(gntNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(gntNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(gntNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(gntNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(gntNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(gntNet_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(gntNet_io_in_1_bits_payload_data),
    .io_in_2_ready(gntNet_io_in_2_ready),
    .io_in_2_valid(gntNet_io_in_2_valid),
    .io_in_2_bits_header_src(gntNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(gntNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(gntNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(gntNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(gntNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(gntNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(gntNet_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(gntNet_io_in_2_bits_payload_data),
    .io_in_3_ready(gntNet_io_in_3_ready),
    .io_in_3_valid(gntNet_io_in_3_valid),
    .io_in_3_bits_header_src(gntNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(gntNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(gntNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(gntNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(gntNet_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(gntNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(gntNet_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(gntNet_io_in_3_bits_payload_data),
    .io_out_0_ready(gntNet_io_out_0_ready),
    .io_out_0_valid(gntNet_io_out_0_valid),
    .io_out_0_bits_header_src(gntNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(gntNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(gntNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_client_xact_id(gntNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_manager_xact_id(gntNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_0_bits_payload_is_builtin_type(gntNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_g_type(gntNet_io_out_0_bits_payload_g_type),
    .io_out_0_bits_payload_data(gntNet_io_out_0_bits_payload_data),
    .io_out_1_ready(gntNet_io_out_1_ready),
    .io_out_1_valid(gntNet_io_out_1_valid),
    .io_out_1_bits_header_src(gntNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(gntNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(gntNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_client_xact_id(gntNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_manager_xact_id(gntNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_1_bits_payload_is_builtin_type(gntNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_g_type(gntNet_io_out_1_bits_payload_g_type),
    .io_out_1_bits_payload_data(gntNet_io_out_1_bits_payload_data),
    .io_out_2_ready(gntNet_io_out_2_ready),
    .io_out_2_valid(gntNet_io_out_2_valid),
    .io_out_2_bits_header_src(gntNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(gntNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(gntNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_client_xact_id(gntNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_manager_xact_id(gntNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_2_bits_payload_is_builtin_type(gntNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_g_type(gntNet_io_out_2_bits_payload_g_type),
    .io_out_2_bits_payload_data(gntNet_io_out_2_bits_payload_data),
    .io_out_3_ready(gntNet_io_out_3_ready),
    .io_out_3_valid(gntNet_io_out_3_valid),
    .io_out_3_bits_header_src(gntNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(gntNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(gntNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_client_xact_id(gntNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_manager_xact_id(gntNet_io_out_3_bits_payload_manager_xact_id),
    .io_out_3_bits_payload_is_builtin_type(gntNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_g_type(gntNet_io_out_3_bits_payload_g_type),
    .io_out_3_bits_payload_data(gntNet_io_out_3_bits_payload_data)
  );
  BasicBus_4 ackNet (
    .clk(ackNet_clk),
    .reset(ackNet_reset),
    .io_in_0_ready(ackNet_io_in_0_ready),
    .io_in_0_valid(ackNet_io_in_0_valid),
    .io_in_0_bits_header_src(ackNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(ackNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(ackNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(ackNet_io_in_1_ready),
    .io_in_1_valid(ackNet_io_in_1_valid),
    .io_in_1_bits_header_src(ackNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(ackNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(ackNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(ackNet_io_in_2_ready),
    .io_in_2_valid(ackNet_io_in_2_valid),
    .io_in_2_bits_header_src(ackNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(ackNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(ackNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(ackNet_io_in_3_ready),
    .io_in_3_valid(ackNet_io_in_3_valid),
    .io_in_3_bits_header_src(ackNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(ackNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(ackNet_io_in_3_bits_payload_manager_xact_id),
    .io_out_0_ready(ackNet_io_out_0_ready),
    .io_out_0_valid(ackNet_io_out_0_valid),
    .io_out_0_bits_header_src(ackNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(ackNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_manager_xact_id(ackNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_1_ready(ackNet_io_out_1_ready),
    .io_out_1_valid(ackNet_io_out_1_valid),
    .io_out_1_bits_header_src(ackNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(ackNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_manager_xact_id(ackNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_2_ready(ackNet_io_out_2_ready),
    .io_out_2_valid(ackNet_io_out_2_valid),
    .io_out_2_bits_header_src(ackNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(ackNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_manager_xact_id(ackNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_3_ready(ackNet_io_out_3_ready),
    .io_out_3_valid(ackNet_io_out_3_valid),
    .io_out_3_bits_header_src(ackNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(ackNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_manager_xact_id(ackNet_io_out_3_bits_payload_manager_xact_id)
  );
  assign io_clients_cached_0_acquire_ready = ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_cached_0_probe_valid = ClientTileLinkNetworkPort_1_io_client_probe_valid;
  assign io_clients_cached_0_probe_bits_addr_block = ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  assign io_clients_cached_0_probe_bits_p_type = ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  assign io_clients_cached_0_release_ready = ClientTileLinkNetworkPort_1_io_client_release_ready;
  assign io_clients_cached_0_grant_valid = ClientTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_cached_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_cached_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_cached_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_cached_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_cached_0_grant_bits_g_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_cached_0_grant_bits_data = ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_clients_cached_0_grant_bits_manager_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id;
  assign io_clients_cached_0_finish_ready = ClientTileLinkNetworkPort_1_io_client_finish_ready;
  assign io_clients_uncached_0_acquire_ready = ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_uncached_0_grant_valid = ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_uncached_0_grant_bits_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_uncached_0_grant_bits_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_uncached_0_grant_bits_manager_xact_id = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_uncached_0_grant_bits_is_builtin_type = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_uncached_0_grant_bits_g_type = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_uncached_0_grant_bits_data = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_2_io_manager_acquire_valid;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_2_io_manager_grant_ready;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_2_io_manager_finish_valid;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_2_io_manager_probe_ready;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_2_io_manager_release_valid;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_2_io_manager_release_bits_data;
  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id;
  assign io_managers_1_acquire_valid = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid;
  assign io_managers_1_acquire_bits_addr_block = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block;
  assign io_managers_1_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id;
  assign io_managers_1_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat;
  assign io_managers_1_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_1_acquire_bits_a_type = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type;
  assign io_managers_1_acquire_bits_union = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union;
  assign io_managers_1_acquire_bits_data = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data;
  assign io_managers_1_acquire_bits_client_id = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id;
  assign io_managers_1_grant_ready = ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready;
  assign io_managers_1_finish_valid = ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid;
  assign io_managers_1_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id;
  assign io_managers_1_probe_ready = ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready;
  assign io_managers_1_release_valid = ManagerTileLinkNetworkPort_1_1_io_manager_release_valid;
  assign io_managers_1_release_bits_addr_beat = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat;
  assign io_managers_1_release_bits_addr_block = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block;
  assign io_managers_1_release_bits_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id;
  assign io_managers_1_release_bits_voluntary = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary;
  assign io_managers_1_release_bits_r_type = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type;
  assign io_managers_1_release_bits_data = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data;
  assign io_managers_1_release_bits_client_id = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id;
  assign TileLinkEnqueuer_4_clk = clk;
  assign TileLinkEnqueuer_4_reset = reset;
  assign TileLinkEnqueuer_4_io_client_acquire_valid = ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_header_src = ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_union = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_data = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_4_io_client_grant_ready = ClientTileLinkNetworkPort_1_io_network_grant_ready;
  assign TileLinkEnqueuer_4_io_client_finish_valid = ClientTileLinkNetworkPort_1_io_network_finish_valid;
  assign TileLinkEnqueuer_4_io_client_finish_bits_header_src = ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_finish_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id = ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_io_client_probe_ready = ClientTileLinkNetworkPort_1_io_network_probe_ready;
  assign TileLinkEnqueuer_4_io_client_release_valid = ClientTileLinkNetworkPort_1_io_network_release_valid;
  assign TileLinkEnqueuer_4_io_client_release_bits_header_src = ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_release_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_r_type = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_data = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_4_io_manager_acquire_ready = T_13624_ready;
  assign TileLinkEnqueuer_4_io_manager_grant_valid = T_17371_valid;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_header_src = T_17371_bits_header_src;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_header_dst = T_17371_bits_header_dst;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat = T_17371_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id = T_17371_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id = T_17371_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type = T_17371_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type = T_17371_bits_payload_g_type;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_data = T_17371_bits_payload_data;
  assign TileLinkEnqueuer_4_io_manager_finish_ready = T_19326_ready;
  assign TileLinkEnqueuer_4_io_manager_probe_valid = T_15939_valid;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_header_src = T_15939_bits_header_src;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_header_dst = T_15939_bits_header_dst;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block = T_15939_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type = T_15939_bits_payload_p_type;
  assign TileLinkEnqueuer_4_io_manager_release_ready = T_15091_ready;
  assign ClientTileLinkNetworkPort_1_clk = clk;
  assign ClientTileLinkNetworkPort_1_reset = reset;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_valid = io_clients_cached_0_acquire_valid;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block = io_clients_cached_0_acquire_bits_addr_block;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id = io_clients_cached_0_acquire_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat = io_clients_cached_0_acquire_bits_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type = io_clients_cached_0_acquire_bits_is_builtin_type;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type = io_clients_cached_0_acquire_bits_a_type;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_union = io_clients_cached_0_acquire_bits_union;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_data = io_clients_cached_0_acquire_bits_data;
  assign ClientTileLinkNetworkPort_1_io_client_probe_ready = io_clients_cached_0_probe_ready;
  assign ClientTileLinkNetworkPort_1_io_client_release_valid = io_clients_cached_0_release_valid;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat = io_clients_cached_0_release_bits_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block = io_clients_cached_0_release_bits_addr_block;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id = io_clients_cached_0_release_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary = io_clients_cached_0_release_bits_voluntary;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_r_type = io_clients_cached_0_release_bits_r_type;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_data = io_clients_cached_0_release_bits_data;
  assign ClientTileLinkNetworkPort_1_io_client_grant_ready = io_clients_cached_0_grant_ready;
  assign ClientTileLinkNetworkPort_1_io_client_finish_valid = io_clients_cached_0_finish_valid;
  assign ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id = io_clients_cached_0_finish_bits_manager_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id = io_clients_cached_0_finish_bits_manager_id;
  assign ClientTileLinkNetworkPort_1_io_network_acquire_ready = TileLinkEnqueuer_4_io_client_acquire_ready;
  assign ClientTileLinkNetworkPort_1_io_network_grant_valid = TileLinkEnqueuer_4_io_client_grant_valid;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src = TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst = TileLinkEnqueuer_4_io_client_grant_bits_header_dst;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data = TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  assign ClientTileLinkNetworkPort_1_io_network_finish_ready = TileLinkEnqueuer_4_io_client_finish_ready;
  assign ClientTileLinkNetworkPort_1_io_network_probe_valid = TileLinkEnqueuer_4_io_client_probe_valid;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src = TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst = TileLinkEnqueuer_4_io_client_probe_bits_header_dst;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  assign ClientTileLinkNetworkPort_1_io_network_release_ready = TileLinkEnqueuer_4_io_client_release_ready;
  assign TileLinkEnqueuer_1_1_clk = clk;
  assign TileLinkEnqueuer_1_1_reset = reset;
  assign TileLinkEnqueuer_1_1_io_client_acquire_valid = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_client_grant_ready = ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready;
  assign TileLinkEnqueuer_1_1_io_client_finish_valid = ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_probe_ready = ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready;
  assign TileLinkEnqueuer_1_1_io_client_release_valid = ClientUncachedTileLinkNetworkPort_1_io_network_release_valid;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_data = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_manager_acquire_ready = T_13794_ready;
  assign TileLinkEnqueuer_1_1_io_manager_grant_valid = T_17936_valid;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src = T_17936_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst = T_17936_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat = T_17936_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id = T_17936_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id = T_17936_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type = T_17936_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type = T_17936_bits_payload_g_type;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data = T_17936_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_manager_finish_ready = T_19466_ready;
  assign TileLinkEnqueuer_1_1_io_manager_probe_valid = T_16484_valid;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src = T_16484_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst = T_16484_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block = T_16484_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type = T_16484_bits_payload_p_type;
  assign TileLinkEnqueuer_1_1_io_manager_release_ready = T_15256_ready;
  assign ClientUncachedTileLinkNetworkPort_1_clk = clk;
  assign ClientUncachedTileLinkNetworkPort_1_reset = reset;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid = io_clients_uncached_0_acquire_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block = io_clients_uncached_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id = io_clients_uncached_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat = io_clients_uncached_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type = io_clients_uncached_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type = io_clients_uncached_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union = io_clients_uncached_0_acquire_bits_union;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data = io_clients_uncached_0_acquire_bits_data;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready = io_clients_uncached_0_grant_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready = TileLinkEnqueuer_1_1_io_client_acquire_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid = TileLinkEnqueuer_1_1_io_client_grant_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src = TileLinkEnqueuer_1_1_io_client_grant_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst = TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready = TileLinkEnqueuer_1_1_io_client_finish_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid = TileLinkEnqueuer_1_1_io_client_probe_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src = TileLinkEnqueuer_1_1_io_client_probe_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst = TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_release_ready = TileLinkEnqueuer_1_1_io_client_release_ready;
  assign ManagerTileLinkNetworkPort_2_clk = clk;
  assign ManagerTileLinkNetworkPort_2_reset = reset;
  assign ManagerTileLinkNetworkPort_2_io_manager_acquire_ready = io_managers_0_acquire_ready;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_valid = io_managers_0_grant_valid;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat = io_managers_0_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id = io_managers_0_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id = io_managers_0_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type = io_managers_0_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type = io_managers_0_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data = io_managers_0_grant_bits_data;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id = io_managers_0_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_finish_ready = io_managers_0_finish_ready;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_valid = io_managers_0_probe_valid;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block = io_managers_0_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type = io_managers_0_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id = io_managers_0_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_release_ready = io_managers_0_release_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_valid = TileLinkEnqueuer_2_1_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src = TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_2_io_network_grant_ready = TileLinkEnqueuer_2_1_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_valid = TileLinkEnqueuer_2_1_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src = TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_probe_ready = TileLinkEnqueuer_2_1_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_release_valid = TileLinkEnqueuer_2_1_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src = TileLinkEnqueuer_2_1_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_2_1_clk = clk;
  assign TileLinkEnqueuer_2_1_reset = reset;
  assign TileLinkEnqueuer_2_1_io_client_acquire_valid = T_12724_valid;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src = T_12724_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst = T_12724_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block = T_12724_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id = T_12724_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat = T_12724_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type = T_12724_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type = T_12724_bits_payload_a_type;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union = T_12724_bits_payload_union;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data = T_12724_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_client_grant_ready = T_16801_ready;
  assign TileLinkEnqueuer_2_1_io_client_finish_valid = T_18486_valid;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_header_src = T_18486_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst = T_18486_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id = T_18486_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_probe_ready = T_15409_ready;
  assign TileLinkEnqueuer_2_1_io_client_release_valid = T_14201_valid;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_header_src = T_14201_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_header_dst = T_14201_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat = T_14201_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block = T_14201_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id = T_14201_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary = T_14201_bits_payload_voluntary;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type = T_14201_bits_payload_r_type;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_data = T_14201_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_manager_acquire_ready = ManagerTileLinkNetworkPort_2_io_network_acquire_ready;
  assign TileLinkEnqueuer_2_1_io_manager_grant_valid = ManagerTileLinkNetworkPort_2_io_network_grant_valid;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_manager_finish_ready = ManagerTileLinkNetworkPort_2_io_network_finish_ready;
  assign TileLinkEnqueuer_2_1_io_manager_probe_valid = ManagerTileLinkNetworkPort_2_io_network_probe_valid;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_2_1_io_manager_release_ready = ManagerTileLinkNetworkPort_2_io_network_release_ready;
  assign ManagerTileLinkNetworkPort_1_1_clk = clk;
  assign ManagerTileLinkNetworkPort_1_1_reset = reset;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready = io_managers_1_acquire_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid = io_managers_1_grant_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat = io_managers_1_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id = io_managers_1_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id = io_managers_1_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type = io_managers_1_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type = io_managers_1_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data = io_managers_1_grant_bits_data;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id = io_managers_1_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready = io_managers_1_finish_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid = io_managers_1_probe_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block = io_managers_1_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type = io_managers_1_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id = io_managers_1_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_release_ready = io_managers_1_release_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid = TileLinkEnqueuer_3_1_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src = TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_1_1_io_network_grant_ready = TileLinkEnqueuer_3_1_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_valid = TileLinkEnqueuer_3_1_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src = TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_probe_ready = TileLinkEnqueuer_3_1_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_valid = TileLinkEnqueuer_3_1_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src = TileLinkEnqueuer_3_1_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_3_1_clk = clk;
  assign TileLinkEnqueuer_3_1_reset = reset;
  assign TileLinkEnqueuer_3_1_io_client_acquire_valid = T_13294_valid;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src = T_13294_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst = T_13294_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block = T_13294_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id = T_13294_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat = T_13294_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type = T_13294_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type = T_13294_bits_payload_a_type;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union = T_13294_bits_payload_union;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data = T_13294_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_client_grant_ready = T_16966_ready;
  assign TileLinkEnqueuer_3_1_io_client_finish_valid = T_19026_valid;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_header_src = T_19026_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst = T_19026_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id = T_19026_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_probe_ready = T_15554_ready;
  assign TileLinkEnqueuer_3_1_io_client_release_valid = T_14766_valid;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_header_src = T_14766_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_header_dst = T_14766_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat = T_14766_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block = T_14766_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id = T_14766_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary = T_14766_bits_payload_voluntary;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type = T_14766_bits_payload_r_type;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_data = T_14766_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_manager_acquire_ready = ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready;
  assign TileLinkEnqueuer_3_1_io_manager_grant_valid = ManagerTileLinkNetworkPort_1_1_io_network_grant_valid;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_manager_finish_ready = ManagerTileLinkNetworkPort_1_1_io_network_finish_ready;
  assign TileLinkEnqueuer_3_1_io_manager_probe_valid = ManagerTileLinkNetworkPort_1_1_io_network_probe_valid;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_3_1_io_manager_release_ready = ManagerTileLinkNetworkPort_1_1_io_network_release_ready;
  assign acqNet_clk = clk;
  assign acqNet_reset = reset;
  assign acqNet_io_in_0_valid = 1'h0;
  assign acqNet_io_in_0_bits_header_src = GEN_0;
  assign acqNet_io_in_0_bits_header_dst = GEN_1;
  assign acqNet_io_in_0_bits_payload_addr_block = GEN_2;
  assign acqNet_io_in_0_bits_payload_client_xact_id = GEN_3;
  assign acqNet_io_in_0_bits_payload_addr_beat = GEN_4;
  assign acqNet_io_in_0_bits_payload_is_builtin_type = GEN_5;
  assign acqNet_io_in_0_bits_payload_a_type = GEN_6;
  assign acqNet_io_in_0_bits_payload_union = GEN_7;
  assign acqNet_io_in_0_bits_payload_data = GEN_8;
  assign acqNet_io_in_1_valid = 1'h0;
  assign acqNet_io_in_1_bits_header_src = GEN_9;
  assign acqNet_io_in_1_bits_header_dst = GEN_10;
  assign acqNet_io_in_1_bits_payload_addr_block = GEN_11;
  assign acqNet_io_in_1_bits_payload_client_xact_id = GEN_12;
  assign acqNet_io_in_1_bits_payload_addr_beat = GEN_13;
  assign acqNet_io_in_1_bits_payload_is_builtin_type = GEN_14;
  assign acqNet_io_in_1_bits_payload_a_type = GEN_15;
  assign acqNet_io_in_1_bits_payload_union = GEN_16;
  assign acqNet_io_in_1_bits_payload_data = GEN_17;
  assign acqNet_io_in_2_valid = T_13624_valid;
  assign acqNet_io_in_2_bits_header_src = T_13624_bits_header_src;
  assign acqNet_io_in_2_bits_header_dst = T_13624_bits_header_dst;
  assign acqNet_io_in_2_bits_payload_addr_block = T_13624_bits_payload_addr_block;
  assign acqNet_io_in_2_bits_payload_client_xact_id = T_13624_bits_payload_client_xact_id;
  assign acqNet_io_in_2_bits_payload_addr_beat = T_13624_bits_payload_addr_beat;
  assign acqNet_io_in_2_bits_payload_is_builtin_type = T_13624_bits_payload_is_builtin_type;
  assign acqNet_io_in_2_bits_payload_a_type = T_13624_bits_payload_a_type;
  assign acqNet_io_in_2_bits_payload_union = T_13624_bits_payload_union;
  assign acqNet_io_in_2_bits_payload_data = T_13624_bits_payload_data;
  assign acqNet_io_in_3_valid = T_13794_valid;
  assign acqNet_io_in_3_bits_header_src = T_13794_bits_header_src;
  assign acqNet_io_in_3_bits_header_dst = T_13794_bits_header_dst;
  assign acqNet_io_in_3_bits_payload_addr_block = T_13794_bits_payload_addr_block;
  assign acqNet_io_in_3_bits_payload_client_xact_id = T_13794_bits_payload_client_xact_id;
  assign acqNet_io_in_3_bits_payload_addr_beat = T_13794_bits_payload_addr_beat;
  assign acqNet_io_in_3_bits_payload_is_builtin_type = T_13794_bits_payload_is_builtin_type;
  assign acqNet_io_in_3_bits_payload_a_type = T_13794_bits_payload_a_type;
  assign acqNet_io_in_3_bits_payload_union = T_13794_bits_payload_union;
  assign acqNet_io_in_3_bits_payload_data = T_13794_bits_payload_data;
  assign acqNet_io_out_0_ready = T_12724_ready;
  assign acqNet_io_out_1_ready = T_13294_ready;
  assign acqNet_io_out_2_ready = 1'h0;
  assign acqNet_io_out_3_ready = 1'h0;
  assign relNet_clk = clk;
  assign relNet_reset = reset;
  assign relNet_io_in_0_valid = 1'h0;
  assign relNet_io_in_0_bits_header_src = GEN_18;
  assign relNet_io_in_0_bits_header_dst = GEN_19;
  assign relNet_io_in_0_bits_payload_addr_beat = GEN_20;
  assign relNet_io_in_0_bits_payload_addr_block = GEN_21;
  assign relNet_io_in_0_bits_payload_client_xact_id = GEN_22;
  assign relNet_io_in_0_bits_payload_voluntary = GEN_23;
  assign relNet_io_in_0_bits_payload_r_type = GEN_24;
  assign relNet_io_in_0_bits_payload_data = GEN_25;
  assign relNet_io_in_1_valid = 1'h0;
  assign relNet_io_in_1_bits_header_src = GEN_26;
  assign relNet_io_in_1_bits_header_dst = GEN_27;
  assign relNet_io_in_1_bits_payload_addr_beat = GEN_28;
  assign relNet_io_in_1_bits_payload_addr_block = GEN_29;
  assign relNet_io_in_1_bits_payload_client_xact_id = GEN_30;
  assign relNet_io_in_1_bits_payload_voluntary = GEN_31;
  assign relNet_io_in_1_bits_payload_r_type = GEN_32;
  assign relNet_io_in_1_bits_payload_data = GEN_33;
  assign relNet_io_in_2_valid = T_15091_valid;
  assign relNet_io_in_2_bits_header_src = T_15091_bits_header_src;
  assign relNet_io_in_2_bits_header_dst = T_15091_bits_header_dst;
  assign relNet_io_in_2_bits_payload_addr_beat = T_15091_bits_payload_addr_beat;
  assign relNet_io_in_2_bits_payload_addr_block = T_15091_bits_payload_addr_block;
  assign relNet_io_in_2_bits_payload_client_xact_id = T_15091_bits_payload_client_xact_id;
  assign relNet_io_in_2_bits_payload_voluntary = T_15091_bits_payload_voluntary;
  assign relNet_io_in_2_bits_payload_r_type = T_15091_bits_payload_r_type;
  assign relNet_io_in_2_bits_payload_data = T_15091_bits_payload_data;
  assign relNet_io_in_3_valid = T_15256_valid;
  assign relNet_io_in_3_bits_header_src = T_15256_bits_header_src;
  assign relNet_io_in_3_bits_header_dst = T_15256_bits_header_dst;
  assign relNet_io_in_3_bits_payload_addr_beat = T_15256_bits_payload_addr_beat;
  assign relNet_io_in_3_bits_payload_addr_block = T_15256_bits_payload_addr_block;
  assign relNet_io_in_3_bits_payload_client_xact_id = T_15256_bits_payload_client_xact_id;
  assign relNet_io_in_3_bits_payload_voluntary = T_15256_bits_payload_voluntary;
  assign relNet_io_in_3_bits_payload_r_type = T_15256_bits_payload_r_type;
  assign relNet_io_in_3_bits_payload_data = T_15256_bits_payload_data;
  assign relNet_io_out_0_ready = T_14201_ready;
  assign relNet_io_out_1_ready = T_14766_ready;
  assign relNet_io_out_2_ready = 1'h0;
  assign relNet_io_out_3_ready = 1'h0;
  assign prbNet_clk = clk;
  assign prbNet_reset = reset;
  assign prbNet_io_in_0_valid = T_15409_valid;
  assign prbNet_io_in_0_bits_header_src = T_15409_bits_header_src;
  assign prbNet_io_in_0_bits_header_dst = T_15409_bits_header_dst;
  assign prbNet_io_in_0_bits_payload_addr_block = T_15409_bits_payload_addr_block;
  assign prbNet_io_in_0_bits_payload_p_type = T_15409_bits_payload_p_type;
  assign prbNet_io_in_1_valid = T_15554_valid;
  assign prbNet_io_in_1_bits_header_src = T_15554_bits_header_src;
  assign prbNet_io_in_1_bits_header_dst = T_15554_bits_header_dst;
  assign prbNet_io_in_1_bits_payload_addr_block = T_15554_bits_payload_addr_block;
  assign prbNet_io_in_1_bits_payload_p_type = T_15554_bits_payload_p_type;
  assign prbNet_io_in_2_valid = 1'h0;
  assign prbNet_io_in_2_bits_header_src = GEN_34;
  assign prbNet_io_in_2_bits_header_dst = GEN_35;
  assign prbNet_io_in_2_bits_payload_addr_block = GEN_36;
  assign prbNet_io_in_2_bits_payload_p_type = GEN_37;
  assign prbNet_io_in_3_valid = 1'h0;
  assign prbNet_io_in_3_bits_header_src = GEN_38;
  assign prbNet_io_in_3_bits_header_dst = GEN_39;
  assign prbNet_io_in_3_bits_payload_addr_block = GEN_40;
  assign prbNet_io_in_3_bits_payload_p_type = GEN_41;
  assign prbNet_io_out_0_ready = 1'h0;
  assign prbNet_io_out_1_ready = 1'h0;
  assign prbNet_io_out_2_ready = T_15939_ready;
  assign prbNet_io_out_3_ready = T_16484_ready;
  assign gntNet_clk = clk;
  assign gntNet_reset = reset;
  assign gntNet_io_in_0_valid = T_16801_valid;
  assign gntNet_io_in_0_bits_header_src = T_16801_bits_header_src;
  assign gntNet_io_in_0_bits_header_dst = T_16801_bits_header_dst;
  assign gntNet_io_in_0_bits_payload_addr_beat = T_16801_bits_payload_addr_beat;
  assign gntNet_io_in_0_bits_payload_client_xact_id = T_16801_bits_payload_client_xact_id;
  assign gntNet_io_in_0_bits_payload_manager_xact_id = T_16801_bits_payload_manager_xact_id;
  assign gntNet_io_in_0_bits_payload_is_builtin_type = T_16801_bits_payload_is_builtin_type;
  assign gntNet_io_in_0_bits_payload_g_type = T_16801_bits_payload_g_type;
  assign gntNet_io_in_0_bits_payload_data = T_16801_bits_payload_data;
  assign gntNet_io_in_1_valid = T_16966_valid;
  assign gntNet_io_in_1_bits_header_src = T_16966_bits_header_src;
  assign gntNet_io_in_1_bits_header_dst = T_16966_bits_header_dst;
  assign gntNet_io_in_1_bits_payload_addr_beat = T_16966_bits_payload_addr_beat;
  assign gntNet_io_in_1_bits_payload_client_xact_id = T_16966_bits_payload_client_xact_id;
  assign gntNet_io_in_1_bits_payload_manager_xact_id = T_16966_bits_payload_manager_xact_id;
  assign gntNet_io_in_1_bits_payload_is_builtin_type = T_16966_bits_payload_is_builtin_type;
  assign gntNet_io_in_1_bits_payload_g_type = T_16966_bits_payload_g_type;
  assign gntNet_io_in_1_bits_payload_data = T_16966_bits_payload_data;
  assign gntNet_io_in_2_valid = 1'h0;
  assign gntNet_io_in_2_bits_header_src = GEN_42;
  assign gntNet_io_in_2_bits_header_dst = GEN_43;
  assign gntNet_io_in_2_bits_payload_addr_beat = GEN_44;
  assign gntNet_io_in_2_bits_payload_client_xact_id = GEN_45;
  assign gntNet_io_in_2_bits_payload_manager_xact_id = GEN_46;
  assign gntNet_io_in_2_bits_payload_is_builtin_type = GEN_47;
  assign gntNet_io_in_2_bits_payload_g_type = GEN_48;
  assign gntNet_io_in_2_bits_payload_data = GEN_49;
  assign gntNet_io_in_3_valid = 1'h0;
  assign gntNet_io_in_3_bits_header_src = GEN_50;
  assign gntNet_io_in_3_bits_header_dst = GEN_51;
  assign gntNet_io_in_3_bits_payload_addr_beat = GEN_52;
  assign gntNet_io_in_3_bits_payload_client_xact_id = GEN_53;
  assign gntNet_io_in_3_bits_payload_manager_xact_id = GEN_54;
  assign gntNet_io_in_3_bits_payload_is_builtin_type = GEN_55;
  assign gntNet_io_in_3_bits_payload_g_type = GEN_56;
  assign gntNet_io_in_3_bits_payload_data = GEN_57;
  assign gntNet_io_out_0_ready = 1'h0;
  assign gntNet_io_out_1_ready = 1'h0;
  assign gntNet_io_out_2_ready = T_17371_ready;
  assign gntNet_io_out_3_ready = T_17936_ready;
  assign ackNet_clk = clk;
  assign ackNet_reset = reset;
  assign ackNet_io_in_0_valid = 1'h0;
  assign ackNet_io_in_0_bits_header_src = GEN_58;
  assign ackNet_io_in_0_bits_header_dst = GEN_59;
  assign ackNet_io_in_0_bits_payload_manager_xact_id = GEN_60;
  assign ackNet_io_in_1_valid = 1'h0;
  assign ackNet_io_in_1_bits_header_src = GEN_61;
  assign ackNet_io_in_1_bits_header_dst = GEN_62;
  assign ackNet_io_in_1_bits_payload_manager_xact_id = GEN_63;
  assign ackNet_io_in_2_valid = T_19326_valid;
  assign ackNet_io_in_2_bits_header_src = T_19326_bits_header_src;
  assign ackNet_io_in_2_bits_header_dst = T_19326_bits_header_dst;
  assign ackNet_io_in_2_bits_payload_manager_xact_id = T_19326_bits_payload_manager_xact_id;
  assign ackNet_io_in_3_valid = T_19466_valid;
  assign ackNet_io_in_3_bits_header_src = T_19466_bits_header_src;
  assign ackNet_io_in_3_bits_header_dst = T_19466_bits_header_dst;
  assign ackNet_io_in_3_bits_payload_manager_xact_id = T_19466_bits_payload_manager_xact_id;
  assign ackNet_io_out_0_ready = T_18486_ready;
  assign ackNet_io_out_1_ready = T_19026_ready;
  assign ackNet_io_out_2_ready = 1'h0;
  assign ackNet_io_out_3_ready = 1'h0;
  assign T_12724_ready = TileLinkEnqueuer_2_1_io_client_acquire_ready;
  assign T_12724_valid = acqNet_io_out_0_valid;
  assign T_12724_bits_header_src = T_12953;
  assign T_12724_bits_header_dst = acqNet_io_out_0_bits_header_dst;
  assign T_12724_bits_payload_addr_block = acqNet_io_out_0_bits_payload_addr_block;
  assign T_12724_bits_payload_client_xact_id = acqNet_io_out_0_bits_payload_client_xact_id;
  assign T_12724_bits_payload_addr_beat = acqNet_io_out_0_bits_payload_addr_beat;
  assign T_12724_bits_payload_is_builtin_type = acqNet_io_out_0_bits_payload_is_builtin_type;
  assign T_12724_bits_payload_a_type = acqNet_io_out_0_bits_payload_a_type;
  assign T_12724_bits_payload_union = acqNet_io_out_0_bits_payload_union;
  assign T_12724_bits_payload_data = acqNet_io_out_0_bits_payload_data;
  assign T_12952 = acqNet_io_out_0_bits_header_src - 2'h2;
  assign T_12953 = T_12952[1:0];
  assign T_13294_ready = TileLinkEnqueuer_3_1_io_client_acquire_ready;
  assign T_13294_valid = acqNet_io_out_1_valid;
  assign T_13294_bits_header_src = T_13523;
  assign T_13294_bits_header_dst = acqNet_io_out_1_bits_header_dst;
  assign T_13294_bits_payload_addr_block = acqNet_io_out_1_bits_payload_addr_block;
  assign T_13294_bits_payload_client_xact_id = acqNet_io_out_1_bits_payload_client_xact_id;
  assign T_13294_bits_payload_addr_beat = acqNet_io_out_1_bits_payload_addr_beat;
  assign T_13294_bits_payload_is_builtin_type = acqNet_io_out_1_bits_payload_is_builtin_type;
  assign T_13294_bits_payload_a_type = acqNet_io_out_1_bits_payload_a_type;
  assign T_13294_bits_payload_union = acqNet_io_out_1_bits_payload_union;
  assign T_13294_bits_payload_data = acqNet_io_out_1_bits_payload_data;
  assign T_13522 = acqNet_io_out_1_bits_header_src - 2'h2;
  assign T_13523 = T_13522[1:0];
  assign T_13624_ready = acqNet_io_in_2_ready;
  assign T_13624_valid = TileLinkEnqueuer_4_io_manager_acquire_valid;
  assign T_13624_bits_header_src = T_13693;
  assign T_13624_bits_header_dst = TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst;
  assign T_13624_bits_payload_addr_block = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block;
  assign T_13624_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id;
  assign T_13624_bits_payload_addr_beat = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat;
  assign T_13624_bits_payload_is_builtin_type = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_13624_bits_payload_a_type = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type;
  assign T_13624_bits_payload_union = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union;
  assign T_13624_bits_payload_data = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data;
  assign T_13692 = TileLinkEnqueuer_4_io_manager_acquire_bits_header_src + 2'h2;
  assign T_13693 = T_13692[1:0];
  assign T_13794_ready = acqNet_io_in_3_ready;
  assign T_13794_valid = TileLinkEnqueuer_1_1_io_manager_acquire_valid;
  assign T_13794_bits_header_src = T_13863;
  assign T_13794_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst;
  assign T_13794_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block;
  assign T_13794_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id;
  assign T_13794_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat;
  assign T_13794_bits_payload_is_builtin_type = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_13794_bits_payload_a_type = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type;
  assign T_13794_bits_payload_union = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union;
  assign T_13794_bits_payload_data = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data;
  assign T_13862 = TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src + 2'h2;
  assign T_13863 = T_13862[1:0];
  assign T_14201_ready = TileLinkEnqueuer_2_1_io_client_release_ready;
  assign T_14201_valid = relNet_io_out_0_valid;
  assign T_14201_bits_header_src = T_14428;
  assign T_14201_bits_header_dst = relNet_io_out_0_bits_header_dst;
  assign T_14201_bits_payload_addr_beat = relNet_io_out_0_bits_payload_addr_beat;
  assign T_14201_bits_payload_addr_block = relNet_io_out_0_bits_payload_addr_block;
  assign T_14201_bits_payload_client_xact_id = relNet_io_out_0_bits_payload_client_xact_id;
  assign T_14201_bits_payload_voluntary = relNet_io_out_0_bits_payload_voluntary;
  assign T_14201_bits_payload_r_type = relNet_io_out_0_bits_payload_r_type;
  assign T_14201_bits_payload_data = relNet_io_out_0_bits_payload_data;
  assign T_14427 = relNet_io_out_0_bits_header_src - 2'h2;
  assign T_14428 = T_14427[1:0];
  assign T_14766_ready = TileLinkEnqueuer_3_1_io_client_release_ready;
  assign T_14766_valid = relNet_io_out_1_valid;
  assign T_14766_bits_header_src = T_14993;
  assign T_14766_bits_header_dst = relNet_io_out_1_bits_header_dst;
  assign T_14766_bits_payload_addr_beat = relNet_io_out_1_bits_payload_addr_beat;
  assign T_14766_bits_payload_addr_block = relNet_io_out_1_bits_payload_addr_block;
  assign T_14766_bits_payload_client_xact_id = relNet_io_out_1_bits_payload_client_xact_id;
  assign T_14766_bits_payload_voluntary = relNet_io_out_1_bits_payload_voluntary;
  assign T_14766_bits_payload_r_type = relNet_io_out_1_bits_payload_r_type;
  assign T_14766_bits_payload_data = relNet_io_out_1_bits_payload_data;
  assign T_14992 = relNet_io_out_1_bits_header_src - 2'h2;
  assign T_14993 = T_14992[1:0];
  assign T_15091_ready = relNet_io_in_2_ready;
  assign T_15091_valid = TileLinkEnqueuer_4_io_manager_release_valid;
  assign T_15091_bits_header_src = T_15158;
  assign T_15091_bits_header_dst = TileLinkEnqueuer_4_io_manager_release_bits_header_dst;
  assign T_15091_bits_payload_addr_beat = TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat;
  assign T_15091_bits_payload_addr_block = TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block;
  assign T_15091_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id;
  assign T_15091_bits_payload_voluntary = TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary;
  assign T_15091_bits_payload_r_type = TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type;
  assign T_15091_bits_payload_data = TileLinkEnqueuer_4_io_manager_release_bits_payload_data;
  assign T_15157 = TileLinkEnqueuer_4_io_manager_release_bits_header_src + 2'h2;
  assign T_15158 = T_15157[1:0];
  assign T_15256_ready = relNet_io_in_3_ready;
  assign T_15256_valid = TileLinkEnqueuer_1_1_io_manager_release_valid;
  assign T_15256_bits_header_src = T_15323;
  assign T_15256_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst;
  assign T_15256_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat;
  assign T_15256_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block;
  assign T_15256_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id;
  assign T_15256_bits_payload_voluntary = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary;
  assign T_15256_bits_payload_r_type = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type;
  assign T_15256_bits_payload_data = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data;
  assign T_15322 = TileLinkEnqueuer_1_1_io_manager_release_bits_header_src + 2'h2;
  assign T_15323 = T_15322[1:0];
  assign T_15409_ready = prbNet_io_in_0_ready;
  assign T_15409_valid = TileLinkEnqueuer_2_1_io_client_probe_valid;
  assign T_15409_bits_header_src = TileLinkEnqueuer_2_1_io_client_probe_bits_header_src;
  assign T_15409_bits_header_dst = T_15468;
  assign T_15409_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block;
  assign T_15409_bits_payload_p_type = TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type;
  assign T_15467 = TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst + 2'h2;
  assign T_15468 = T_15467[1:0];
  assign T_15554_ready = prbNet_io_in_1_ready;
  assign T_15554_valid = TileLinkEnqueuer_3_1_io_client_probe_valid;
  assign T_15554_bits_header_src = TileLinkEnqueuer_3_1_io_client_probe_bits_header_src;
  assign T_15554_bits_header_dst = T_15613;
  assign T_15554_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block;
  assign T_15554_bits_payload_p_type = TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type;
  assign T_15612 = TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst + 2'h2;
  assign T_15613 = T_15612[1:0];
  assign T_15939_ready = TileLinkEnqueuer_4_io_manager_probe_ready;
  assign T_15939_valid = prbNet_io_out_2_valid;
  assign T_15939_bits_header_src = prbNet_io_out_2_bits_header_src;
  assign T_15939_bits_header_dst = T_16158;
  assign T_15939_bits_payload_addr_block = prbNet_io_out_2_bits_payload_addr_block;
  assign T_15939_bits_payload_p_type = prbNet_io_out_2_bits_payload_p_type;
  assign T_16157 = prbNet_io_out_2_bits_header_dst - 2'h2;
  assign T_16158 = T_16157[1:0];
  assign T_16484_ready = TileLinkEnqueuer_1_1_io_manager_probe_ready;
  assign T_16484_valid = prbNet_io_out_3_valid;
  assign T_16484_bits_header_src = prbNet_io_out_3_bits_header_src;
  assign T_16484_bits_header_dst = T_16703;
  assign T_16484_bits_payload_addr_block = prbNet_io_out_3_bits_payload_addr_block;
  assign T_16484_bits_payload_p_type = prbNet_io_out_3_bits_payload_p_type;
  assign T_16702 = prbNet_io_out_3_bits_header_dst - 2'h2;
  assign T_16703 = T_16702[1:0];
  assign T_16801_ready = gntNet_io_in_0_ready;
  assign T_16801_valid = TileLinkEnqueuer_2_1_io_client_grant_valid;
  assign T_16801_bits_header_src = TileLinkEnqueuer_2_1_io_client_grant_bits_header_src;
  assign T_16801_bits_header_dst = T_16868;
  assign T_16801_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat;
  assign T_16801_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id;
  assign T_16801_bits_payload_manager_xact_id = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id;
  assign T_16801_bits_payload_is_builtin_type = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type;
  assign T_16801_bits_payload_g_type = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type;
  assign T_16801_bits_payload_data = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data;
  assign T_16867 = TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst + 2'h2;
  assign T_16868 = T_16867[1:0];
  assign T_16966_ready = gntNet_io_in_1_ready;
  assign T_16966_valid = TileLinkEnqueuer_3_1_io_client_grant_valid;
  assign T_16966_bits_header_src = TileLinkEnqueuer_3_1_io_client_grant_bits_header_src;
  assign T_16966_bits_header_dst = T_17033;
  assign T_16966_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat;
  assign T_16966_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id;
  assign T_16966_bits_payload_manager_xact_id = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id;
  assign T_16966_bits_payload_is_builtin_type = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type;
  assign T_16966_bits_payload_g_type = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type;
  assign T_16966_bits_payload_data = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data;
  assign T_17032 = TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst + 2'h2;
  assign T_17033 = T_17032[1:0];
  assign T_17371_ready = TileLinkEnqueuer_4_io_manager_grant_ready;
  assign T_17371_valid = gntNet_io_out_2_valid;
  assign T_17371_bits_header_src = gntNet_io_out_2_bits_header_src;
  assign T_17371_bits_header_dst = T_17598;
  assign T_17371_bits_payload_addr_beat = gntNet_io_out_2_bits_payload_addr_beat;
  assign T_17371_bits_payload_client_xact_id = gntNet_io_out_2_bits_payload_client_xact_id;
  assign T_17371_bits_payload_manager_xact_id = gntNet_io_out_2_bits_payload_manager_xact_id;
  assign T_17371_bits_payload_is_builtin_type = gntNet_io_out_2_bits_payload_is_builtin_type;
  assign T_17371_bits_payload_g_type = gntNet_io_out_2_bits_payload_g_type;
  assign T_17371_bits_payload_data = gntNet_io_out_2_bits_payload_data;
  assign T_17597 = gntNet_io_out_2_bits_header_dst - 2'h2;
  assign T_17598 = T_17597[1:0];
  assign T_17936_ready = TileLinkEnqueuer_1_1_io_manager_grant_ready;
  assign T_17936_valid = gntNet_io_out_3_valid;
  assign T_17936_bits_header_src = gntNet_io_out_3_bits_header_src;
  assign T_17936_bits_header_dst = T_18163;
  assign T_17936_bits_payload_addr_beat = gntNet_io_out_3_bits_payload_addr_beat;
  assign T_17936_bits_payload_client_xact_id = gntNet_io_out_3_bits_payload_client_xact_id;
  assign T_17936_bits_payload_manager_xact_id = gntNet_io_out_3_bits_payload_manager_xact_id;
  assign T_17936_bits_payload_is_builtin_type = gntNet_io_out_3_bits_payload_is_builtin_type;
  assign T_17936_bits_payload_g_type = gntNet_io_out_3_bits_payload_g_type;
  assign T_17936_bits_payload_data = gntNet_io_out_3_bits_payload_data;
  assign T_18162 = gntNet_io_out_3_bits_header_dst - 2'h2;
  assign T_18163 = T_18162[1:0];
  assign T_18486_ready = TileLinkEnqueuer_2_1_io_client_finish_ready;
  assign T_18486_valid = ackNet_io_out_0_valid;
  assign T_18486_bits_header_src = T_18703;
  assign T_18486_bits_header_dst = ackNet_io_out_0_bits_header_dst;
  assign T_18486_bits_payload_manager_xact_id = ackNet_io_out_0_bits_payload_manager_xact_id;
  assign T_18702 = ackNet_io_out_0_bits_header_src - 2'h2;
  assign T_18703 = T_18702[1:0];
  assign T_19026_ready = TileLinkEnqueuer_3_1_io_client_finish_ready;
  assign T_19026_valid = ackNet_io_out_1_valid;
  assign T_19026_bits_header_src = T_19243;
  assign T_19026_bits_header_dst = ackNet_io_out_1_bits_header_dst;
  assign T_19026_bits_payload_manager_xact_id = ackNet_io_out_1_bits_payload_manager_xact_id;
  assign T_19242 = ackNet_io_out_1_bits_header_src - 2'h2;
  assign T_19243 = T_19242[1:0];
  assign T_19326_ready = ackNet_io_in_2_ready;
  assign T_19326_valid = TileLinkEnqueuer_4_io_manager_finish_valid;
  assign T_19326_bits_header_src = T_19383;
  assign T_19326_bits_header_dst = TileLinkEnqueuer_4_io_manager_finish_bits_header_dst;
  assign T_19326_bits_payload_manager_xact_id = TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id;
  assign T_19382 = TileLinkEnqueuer_4_io_manager_finish_bits_header_src + 2'h2;
  assign T_19383 = T_19382[1:0];
  assign T_19466_ready = ackNet_io_in_3_ready;
  assign T_19466_valid = TileLinkEnqueuer_1_1_io_manager_finish_valid;
  assign T_19466_bits_header_src = T_19523;
  assign T_19466_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst;
  assign T_19466_bits_payload_manager_xact_id = TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id;
  assign T_19522 = TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src + 2'h2;
  assign T_19523 = T_19522[1:0];
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_0 = GEN_64[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_65[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_66[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_67[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_4 = GEN_68[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_5 = GEN_69[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_6 = GEN_70[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_7 = GEN_71[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_8 = GEN_72[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_9 = GEN_73[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_10 = GEN_74[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_11 = GEN_75[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_12 = GEN_76[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_13 = GEN_77[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_14 = GEN_78[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_15 = GEN_79[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_16 = GEN_80[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_17 = GEN_81[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_18 = GEN_82[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_19 = GEN_83[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_20 = GEN_84[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_21 = GEN_85[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_22 = GEN_86[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_23 = GEN_87[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_24 = GEN_88[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_25 = GEN_89[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_26 = GEN_90[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_27 = GEN_91[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_28 = GEN_92[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_29 = GEN_93[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_94[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_95[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_32 = GEN_96[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_33 = GEN_97[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_34 = GEN_98[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_35 = GEN_99[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_36 = GEN_100[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_37 = GEN_101[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_38 = GEN_102[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_39 = GEN_103[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_40 = GEN_104[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_41 = GEN_105[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_42 = GEN_106[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_43 = GEN_107[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_44 = GEN_108[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_45 = GEN_109[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_46 = GEN_110[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_47 = GEN_111[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_48 = GEN_112[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_49 = GEN_113[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_50 = GEN_114[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_51 = GEN_115[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_52 = GEN_116[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_53 = GEN_117[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_54 = GEN_118[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_55 = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_56 = GEN_120[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_57 = GEN_121[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_58 = GEN_122[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_59 = GEN_123[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_60 = GEN_124[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_61 = GEN_125[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_62 = GEN_126[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_63 = GEN_127[1:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_64 = {1{$random}};
  GEN_65 = {1{$random}};
  GEN_66 = {1{$random}};
  GEN_67 = {1{$random}};
  GEN_68 = {1{$random}};
  GEN_69 = {1{$random}};
  GEN_70 = {1{$random}};
  GEN_71 = {1{$random}};
  GEN_72 = {2{$random}};
  GEN_73 = {1{$random}};
  GEN_74 = {1{$random}};
  GEN_75 = {1{$random}};
  GEN_76 = {1{$random}};
  GEN_77 = {1{$random}};
  GEN_78 = {1{$random}};
  GEN_79 = {1{$random}};
  GEN_80 = {1{$random}};
  GEN_81 = {2{$random}};
  GEN_82 = {1{$random}};
  GEN_83 = {1{$random}};
  GEN_84 = {1{$random}};
  GEN_85 = {1{$random}};
  GEN_86 = {1{$random}};
  GEN_87 = {1{$random}};
  GEN_88 = {1{$random}};
  GEN_89 = {2{$random}};
  GEN_90 = {1{$random}};
  GEN_91 = {1{$random}};
  GEN_92 = {1{$random}};
  GEN_93 = {1{$random}};
  GEN_94 = {1{$random}};
  GEN_95 = {1{$random}};
  GEN_96 = {1{$random}};
  GEN_97 = {2{$random}};
  GEN_98 = {1{$random}};
  GEN_99 = {1{$random}};
  GEN_100 = {1{$random}};
  GEN_101 = {1{$random}};
  GEN_102 = {1{$random}};
  GEN_103 = {1{$random}};
  GEN_104 = {1{$random}};
  GEN_105 = {1{$random}};
  GEN_106 = {1{$random}};
  GEN_107 = {1{$random}};
  GEN_108 = {1{$random}};
  GEN_109 = {1{$random}};
  GEN_110 = {1{$random}};
  GEN_111 = {1{$random}};
  GEN_112 = {1{$random}};
  GEN_113 = {2{$random}};
  GEN_114 = {1{$random}};
  GEN_115 = {1{$random}};
  GEN_116 = {1{$random}};
  GEN_117 = {1{$random}};
  GEN_118 = {1{$random}};
  GEN_119 = {1{$random}};
  GEN_120 = {1{$random}};
  GEN_121 = {2{$random}};
  GEN_122 = {1{$random}};
  GEN_123 = {1{$random}};
  GEN_124 = {1{$random}};
  GEN_125 = {1{$random}};
  GEN_126 = {1{$random}};
  GEN_127 = {1{$random}};
  end
`endif
endmodule
module BufferedBroadcastVoluntaryReleaseTracker(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input   io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output  io_inner_grant_bits_client_xact_id,
  output [1:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [1:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input   io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [1:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should,
  output  io_alloc_idle,
  output [25:0] io_alloc_addr_block
);
  wire  all_pending_done;
  reg [3:0] state;
  reg [31:0] GEN_69;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_70;
  reg [2:0] xact_vol_ir_r_type;
  reg [31:0] GEN_71;
  reg  xact_vol_ir_src;
  reg [31:0] GEN_72;
  reg  xact_vol_ir_client_xact_id;
  reg [31:0] GEN_73;
  reg [7:0] pending_irel_data;
  reg [31:0] GEN_74;
  wire  vol_ignt_counter_pending;
  wire [2:0] vol_ignt_counter_up_idx;
  wire  vol_ignt_counter_up_done;
  wire [2:0] vol_ignt_counter_down_idx;
  wire  vol_ignt_counter_down_done;
  reg  pending_orel_send;
  reg [31:0] GEN_75;
  reg [7:0] pending_orel_data;
  reg [31:0] GEN_76;
  wire  vol_ognt_counter_pending;
  wire [2:0] vol_ognt_counter_up_idx;
  wire  vol_ognt_counter_up_done;
  wire [2:0] vol_ognt_counter_down_idx;
  wire  vol_ognt_counter_down_done;
  wire  T_78;
  wire  T_79;
  wire  scoreboard_2;
  reg  sending_orel;
  reg [31:0] GEN_77;
  wire  T_103_sharers;
  wire [1:0] T_149_state;
  wire  coh_inner_sharers;
  wire [1:0] coh_outer_state;
  wire  T_1519;
  wire  T_1520;
  wire  T_1521;
  wire  T_1522;
  wire  T_1524;
  wire  T_1525;
  wire  T_1527;
  wire  T_1528;
  wire  T_1530;
  wire [63:0] T_1544_0;
  wire [63:0] T_1544_1;
  wire [63:0] T_1544_2;
  wire [63:0] T_1544_3;
  wire [63:0] T_1544_4;
  wire [63:0] T_1544_5;
  wire [63:0] T_1544_6;
  wire [63:0] T_1544_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_78;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_79;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_80;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_81;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_82;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_83;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_84;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_85;
  wire  T_1552;
  wire  T_1553;
  wire  T_1554;
  wire  T_1556;
  wire  T_1557;
  wire  T_1559;
  wire  T_1560;
  wire  T_1568;
  wire  T_1572;
  wire  T_1573;
  wire  T_1578;
  wire  T_1580;
  wire  T_1581;
  wire  T_1582;
  wire  T_1583;
  wire  T_1584;
  wire  T_1586;
  reg [2:0] T_1588;
  reg [31:0] GEN_86;
  wire  T_1590;
  wire [3:0] T_1592;
  wire [2:0] T_1593;
  wire [2:0] GEN_2;
  wire  T_1594;
  wire [2:0] T_1595;
  wire  T_1596;
  wire  T_1597;
  wire  T_1600;
  wire  T_1601;
  wire  T_1602;
  wire  T_1603;
  wire [2:0] T_1611_0;
  wire [3:0] GEN_57;
  wire  T_1613;
  wire  T_1615;
  wire  T_1617;
  reg [2:0] T_1619;
  reg [31:0] GEN_87;
  wire  T_1621;
  wire [3:0] T_1623;
  wire [2:0] T_1624;
  wire [2:0] GEN_3;
  wire  T_1625;
  wire [2:0] T_1626;
  wire  T_1627;
  reg  T_1629;
  reg [31:0] GEN_88;
  wire  T_1631;
  wire  T_1632;
  wire [1:0] T_1634;
  wire  T_1635;
  wire  GEN_4;
  wire  T_1637;
  wire  T_1638;
  wire [1:0] T_1640;
  wire  T_1641;
  wire  GEN_5;
  wire  T_1643;
  wire  T_1645;
  wire  T_1646;
  wire [25:0] GEN_6;
  wire [7:0] GEN_7;
  wire [3:0] GEN_8;
  wire  T_1654;
  wire  T_1656;
  wire  T_1657;
  wire  T_1659;
  wire  T_1660;
  wire  T_1661;
  wire  T_1670;
  wire  T_1672;
  wire  T_1673;
  wire [2:0] GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  T_1687;
  wire [7:0] T_1691;
  wire [7:0] T_1692;
  wire [7:0] T_1694;
  wire [7:0] T_1695;
  wire [7:0] T_1696;
  wire [7:0] T_1698;
  wire [2:0] GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [7:0] GEN_15;
  wire  T_1700;
  wire [7:0] T_1717;
  wire [7:0] GEN_16;
  wire [2:0] GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire [7:0] GEN_20;
  wire  T_1718;
  wire  T_1719;
  wire  T_1720;
  wire  T_1721;
  wire  T_1722;
  wire  T_1723;
  wire  T_1724;
  wire  T_1725;
  wire  T_1728;
  wire  T_1730;
  wire  T_1731;
  wire [2:0] T_1763_addr_beat;
  wire [25:0] T_1763_addr_block;
  wire  T_1763_client_xact_id;
  wire  T_1763_voluntary;
  wire [2:0] T_1763_r_type;
  wire [63:0] T_1763_data;
  wire  T_1763_client_id;
  wire [2:0] T_1824_addr_beat;
  wire  T_1824_client_xact_id;
  wire [1:0] T_1824_manager_xact_id;
  wire  T_1824_is_builtin_type;
  wire [3:0] T_1824_g_type;
  wire [63:0] T_1824_data;
  wire  T_1824_client_id;
  wire  T_1861;
  wire [63:0] GEN_0;
  wire [63:0] GEN_21;
  wire [63:0] GEN_22;
  wire [63:0] GEN_23;
  wire [63:0] GEN_24;
  wire [63:0] GEN_25;
  wire [63:0] GEN_26;
  wire [63:0] GEN_27;
  wire [63:0] GEN_28;
  wire [63:0] GEN_30;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  wire [63:0] GEN_36;
  wire [63:0] GEN_37;
  wire [1:0] T_1893_state;
  wire  T_1922;
  wire [7:0] T_1938;
  wire [7:0] T_1939;
  wire  T_1941;
  wire  T_1942;
  wire  T_1943;
  wire  T_1944;
  wire  T_1945;
  wire  T_1946;
  wire  T_1947;
  wire [7:0] T_1951;
  wire [7:0] T_1952;
  wire [7:0] T_1954;
  wire [7:0] T_1955;
  wire [7:0] T_1956;
  wire [7:0] T_1957;
  wire [7:0] GEN_38;
  wire  GEN_39;
  wire  T_1968;
  wire  T_1970;
  wire  T_1971;
  wire  GEN_40;
  wire  T_1983;
  wire  T_1984;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  T_1993;
  wire  T_2001;
  reg [2:0] T_2003;
  reg [31:0] GEN_89;
  wire  T_2005;
  wire [3:0] T_2007;
  wire [2:0] T_2008;
  wire [2:0] GEN_44;
  wire  T_2009;
  wire [2:0] T_2010;
  wire  T_2011;
  wire  T_2012;
  wire  T_2014;
  wire  T_2015;
  wire  T_2016;
  wire [2:0] T_2024_0;
  wire [3:0] GEN_58;
  wire  T_2026;
  wire  T_2028;
  wire  T_2030;
  reg [2:0] T_2032;
  reg [31:0] GEN_90;
  wire  T_2034;
  wire [3:0] T_2036;
  wire [2:0] T_2037;
  wire [2:0] GEN_45;
  wire  T_2038;
  wire [2:0] T_2039;
  wire  T_2040;
  reg  T_2042;
  reg [31:0] GEN_91;
  wire  T_2044;
  wire  T_2045;
  wire [1:0] T_2047;
  wire  T_2048;
  wire  GEN_46;
  wire  T_2050;
  wire  T_2051;
  wire [1:0] T_2053;
  wire  T_2054;
  wire  GEN_47;
  wire  T_2056;
  wire [7:0] T_2065;
  wire  T_2066;
  wire  T_2067;
  wire  T_2068;
  wire  T_2082;
  wire [2:0] T_2083;
  wire [2:0] T_2119_addr_beat;
  wire [25:0] T_2119_addr_block;
  wire [1:0] T_2119_client_xact_id;
  wire  T_2119_voluntary;
  wire [2:0] T_2119_r_type;
  wire [63:0] T_2119_data;
  wire [63:0] GEN_1;
  wire [63:0] GEN_48;
  wire [63:0] GEN_49;
  wire [63:0] GEN_50;
  wire [63:0] GEN_51;
  wire [63:0] GEN_52;
  wire [63:0] GEN_53;
  wire [63:0] GEN_54;
  wire  T_2149;
  wire  T_2150;
  wire  T_2151;
  wire  T_2153;
  wire  T_2155;
  wire [3:0] GEN_56;
  wire [25:0] GEN_29;
  reg [31:0] GEN_92;
  wire [1:0] GEN_55;
  reg [31:0] GEN_93;
  wire  GEN_59;
  reg [31:0] GEN_94;
  wire [25:0] GEN_60;
  reg [31:0] GEN_95;
  wire [1:0] GEN_61;
  reg [31:0] GEN_96;
  wire [2:0] GEN_62;
  reg [31:0] GEN_97;
  wire  GEN_63;
  reg [31:0] GEN_98;
  wire [2:0] GEN_64;
  reg [31:0] GEN_99;
  wire [10:0] GEN_65;
  reg [31:0] GEN_100;
  wire [63:0] GEN_66;
  reg [63:0] GEN_101;
  wire  GEN_67;
  reg [31:0] GEN_102;
  wire  GEN_68;
  reg [31:0] GEN_103;
  assign io_inner_acquire_ready = 1'h0;
  assign io_inner_grant_valid = T_1731;
  assign io_inner_grant_bits_addr_beat = T_1824_addr_beat;
  assign io_inner_grant_bits_client_xact_id = T_1824_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = T_1824_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = T_1824_is_builtin_type;
  assign io_inner_grant_bits_g_type = T_1824_g_type;
  assign io_inner_grant_bits_data = T_1824_data;
  assign io_inner_grant_bits_client_id = T_1824_client_id;
  assign io_inner_finish_ready = 1'h0;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_29;
  assign io_inner_probe_bits_p_type = GEN_55;
  assign io_inner_probe_bits_client_id = GEN_59;
  assign io_inner_release_ready = T_1861;
  assign io_outer_acquire_valid = 1'h0;
  assign io_outer_acquire_bits_addr_block = GEN_60;
  assign io_outer_acquire_bits_client_xact_id = GEN_61;
  assign io_outer_acquire_bits_addr_beat = GEN_62;
  assign io_outer_acquire_bits_is_builtin_type = GEN_63;
  assign io_outer_acquire_bits_a_type = GEN_64;
  assign io_outer_acquire_bits_union = GEN_65;
  assign io_outer_acquire_bits_data = GEN_66;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2068;
  assign io_outer_release_bits_addr_beat = T_2119_addr_beat;
  assign io_outer_release_bits_addr_block = T_2119_addr_block;
  assign io_outer_release_bits_client_xact_id = T_2119_client_xact_id;
  assign io_outer_release_bits_voluntary = T_2119_voluntary;
  assign io_outer_release_bits_r_type = T_2119_r_type;
  assign io_outer_release_bits_data = T_2119_data;
  assign io_outer_grant_ready = vol_ognt_counter_pending;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_67;
  assign io_outer_finish_bits_manager_id = GEN_68;
  assign io_alloc_iacq_matches = T_1554;
  assign io_alloc_iacq_can = 1'h0;
  assign io_alloc_irel_matches = T_1557;
  assign io_alloc_irel_can = T_1519;
  assign io_alloc_oprb_matches = T_1560;
  assign io_alloc_oprb_can = 1'h0;
  assign io_alloc_idle = T_1519;
  assign io_alloc_addr_block = xact_addr_block;
  assign all_pending_done = T_2153;
  assign vol_ignt_counter_pending = T_1643;
  assign vol_ignt_counter_up_idx = T_1595;
  assign vol_ignt_counter_up_done = T_1596;
  assign vol_ignt_counter_down_idx = T_1626;
  assign vol_ignt_counter_down_done = T_1627;
  assign vol_ognt_counter_pending = T_2056;
  assign vol_ognt_counter_up_idx = T_2010;
  assign vol_ognt_counter_up_done = T_2011;
  assign vol_ognt_counter_down_idx = T_2039;
  assign vol_ognt_counter_down_done = T_2040;
  assign T_78 = pending_orel_data != 8'h0;
  assign T_79 = pending_orel_send | T_78;
  assign scoreboard_2 = T_79 | vol_ognt_counter_pending;
  assign T_103_sharers = 1'h0;
  assign T_149_state = 2'h0;
  assign coh_inner_sharers = T_103_sharers;
  assign coh_outer_state = T_149_state;
  assign T_1519 = state == 4'h0;
  assign T_1520 = io_inner_release_ready & io_inner_release_valid;
  assign T_1521 = T_1519 & T_1520;
  assign T_1522 = T_1521 & io_alloc_irel_should;
  assign T_1524 = io_inner_release_bits_voluntary == 1'h0;
  assign T_1525 = T_1522 & T_1524;
  assign T_1527 = T_1525 == 1'h0;
  assign T_1528 = T_1527 | reset;
  assign T_1530 = T_1528 == 1'h0;
  assign T_1544_0 = 64'h0;
  assign T_1544_1 = 64'h0;
  assign T_1544_2 = 64'h0;
  assign T_1544_3 = 64'h0;
  assign T_1544_4 = 64'h0;
  assign T_1544_5 = 64'h0;
  assign T_1544_6 = 64'h0;
  assign T_1544_7 = 64'h0;
  assign T_1552 = state != 4'h0;
  assign T_1553 = io_inner_acquire_bits_addr_block == xact_addr_block;
  assign T_1554 = T_1552 & T_1553;
  assign T_1556 = io_inner_release_bits_addr_block == xact_addr_block;
  assign T_1557 = T_1552 & T_1556;
  assign T_1559 = io_outer_probe_bits_addr_block == xact_addr_block;
  assign T_1560 = T_1552 & T_1559;
  assign T_1568 = scoreboard_2 | vol_ognt_counter_pending;
  assign T_1572 = T_1519 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_1573 = T_1572 & io_inner_release_bits_voluntary;
  assign T_1578 = T_1520 & T_1573;
  assign T_1580 = io_inner_release_bits_r_type == 3'h0;
  assign T_1581 = io_inner_release_bits_r_type == 3'h1;
  assign T_1582 = io_inner_release_bits_r_type == 3'h2;
  assign T_1583 = T_1580 | T_1581;
  assign T_1584 = T_1583 | T_1582;
  assign T_1586 = T_1578 & T_1584;
  assign T_1590 = T_1588 == 3'h7;
  assign T_1592 = T_1588 + 3'h1;
  assign T_1593 = T_1592[2:0];
  assign GEN_2 = T_1586 ? T_1593 : T_1588;
  assign T_1594 = T_1586 & T_1590;
  assign T_1595 = T_1584 ? T_1588 : 3'h0;
  assign T_1596 = T_1584 ? T_1594 : T_1578;
  assign T_1597 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_1600 = io_inner_grant_bits_g_type == 4'h0;
  assign T_1601 = io_inner_grant_bits_is_builtin_type & T_1600;
  assign T_1602 = T_1552 & T_1601;
  assign T_1603 = T_1597 & T_1602;
  assign T_1611_0 = 3'h5;
  assign GEN_57 = {{1'd0}, T_1611_0};
  assign T_1613 = io_inner_grant_bits_g_type == GEN_57;
  assign T_1615 = io_inner_grant_bits_is_builtin_type ? T_1613 : T_1600;
  assign T_1617 = T_1603 & T_1615;
  assign T_1621 = T_1619 == 3'h7;
  assign T_1623 = T_1619 + 3'h1;
  assign T_1624 = T_1623[2:0];
  assign GEN_3 = T_1617 ? T_1624 : T_1619;
  assign T_1625 = T_1617 & T_1621;
  assign T_1626 = T_1615 ? T_1619 : 3'h0;
  assign T_1627 = T_1615 ? T_1625 : T_1603;
  assign T_1631 = T_1627 == 1'h0;
  assign T_1632 = T_1596 & T_1631;
  assign T_1634 = T_1629 + 1'h1;
  assign T_1635 = T_1634[0:0];
  assign GEN_4 = T_1632 ? T_1635 : T_1629;
  assign T_1637 = T_1596 == 1'h0;
  assign T_1638 = T_1627 & T_1637;
  assign T_1640 = T_1629 - 1'h1;
  assign T_1641 = T_1640[0:0];
  assign GEN_5 = T_1638 ? T_1641 : GEN_4;
  assign T_1643 = T_1629 > 1'h0;
  assign T_1645 = T_1519 & io_alloc_irel_should;
  assign T_1646 = T_1645 & io_inner_release_valid;
  assign GEN_6 = T_1646 ? io_inner_release_bits_addr_block : xact_addr_block;
  assign GEN_7 = T_1646 ? 8'hff : pending_irel_data;
  assign GEN_8 = T_1646 ? 4'h7 : state;
  assign T_1654 = T_1556 & io_inner_release_bits_voluntary;
  assign T_1656 = pending_irel_data != 8'h0;
  assign T_1657 = T_1654 & T_1656;
  assign T_1659 = T_1657 & io_inner_release_valid;
  assign T_1660 = T_1646 | T_1659;
  assign T_1661 = T_1660 & io_inner_release_ready;
  assign T_1670 = T_1584 == 1'h0;
  assign T_1672 = io_inner_release_bits_addr_beat == 3'h0;
  assign T_1673 = T_1670 | T_1672;
  assign GEN_9 = io_inner_release_bits_voluntary ? io_inner_release_bits_r_type : xact_vol_ir_r_type;
  assign GEN_10 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_id : xact_vol_ir_src;
  assign GEN_11 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_xact_id : xact_vol_ir_client_xact_id;
  assign T_1687 = T_1520 & T_1584;
  assign T_1691 = T_1687 ? 8'hff : 8'h0;
  assign T_1692 = ~ T_1691;
  assign T_1694 = 8'h1 << io_inner_release_bits_addr_beat;
  assign T_1695 = ~ T_1694;
  assign T_1696 = T_1692 | T_1695;
  assign T_1698 = T_1584 ? T_1696 : 8'h0;
  assign GEN_12 = T_1673 ? GEN_9 : xact_vol_ir_r_type;
  assign GEN_13 = T_1673 ? GEN_10 : xact_vol_ir_src;
  assign GEN_14 = T_1673 ? GEN_11 : xact_vol_ir_client_xact_id;
  assign GEN_15 = T_1673 ? T_1698 : GEN_7;
  assign T_1700 = T_1673 == 1'h0;
  assign T_1717 = pending_irel_data & T_1696;
  assign GEN_16 = T_1700 ? T_1717 : GEN_15;
  assign GEN_17 = T_1661 ? GEN_12 : xact_vol_ir_r_type;
  assign GEN_18 = T_1661 ? GEN_13 : xact_vol_ir_src;
  assign GEN_19 = T_1661 ? GEN_14 : xact_vol_ir_client_xact_id;
  assign GEN_20 = T_1661 ? GEN_16 : GEN_7;
  assign T_1718 = state == 4'h3;
  assign T_1719 = state == 4'h4;
  assign T_1720 = state == 4'h5;
  assign T_1721 = state == 4'h7;
  assign T_1722 = T_1718 | T_1719;
  assign T_1723 = T_1722 | T_1720;
  assign T_1724 = T_1723 | T_1721;
  assign T_1725 = T_1724 & vol_ignt_counter_pending;
  assign T_1728 = T_1656 | T_1568;
  assign T_1730 = T_1728 == 1'h0;
  assign T_1731 = T_1725 & T_1730;
  assign T_1763_addr_beat = 3'h0;
  assign T_1763_addr_block = xact_addr_block;
  assign T_1763_client_xact_id = xact_vol_ir_client_xact_id;
  assign T_1763_voluntary = 1'h1;
  assign T_1763_r_type = xact_vol_ir_r_type;
  assign T_1763_data = 64'h0;
  assign T_1763_client_id = xact_vol_ir_src;
  assign T_1824_addr_beat = 3'h0;
  assign T_1824_client_xact_id = T_1763_client_xact_id;
  assign T_1824_manager_xact_id = 2'h0;
  assign T_1824_is_builtin_type = 1'h1;
  assign T_1824_g_type = 4'h0;
  assign T_1824_data = 64'h0;
  assign T_1824_client_id = T_1763_client_id;
  assign T_1861 = T_1519 | T_1657;
  assign GEN_0 = io_inner_release_bits_data;
  assign GEN_21 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_0;
  assign GEN_22 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_1;
  assign GEN_23 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_2;
  assign GEN_24 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_3;
  assign GEN_25 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_4;
  assign GEN_26 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_5;
  assign GEN_27 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_6;
  assign GEN_28 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_7;
  assign GEN_30 = T_1520 ? GEN_21 : data_buffer_0;
  assign GEN_31 = T_1520 ? GEN_22 : data_buffer_1;
  assign GEN_32 = T_1520 ? GEN_23 : data_buffer_2;
  assign GEN_33 = T_1520 ? GEN_24 : data_buffer_3;
  assign GEN_34 = T_1520 ? GEN_25 : data_buffer_4;
  assign GEN_35 = T_1520 ? GEN_26 : data_buffer_5;
  assign GEN_36 = T_1520 ? GEN_27 : data_buffer_6;
  assign GEN_37 = T_1520 ? GEN_28 : data_buffer_7;
  assign T_1893_state = 2'h2;
  assign T_1922 = T_1552 | io_alloc_irel_should;
  assign T_1938 = T_1691 & T_1694;
  assign T_1939 = pending_orel_data | T_1938;
  assign T_1941 = io_outer_release_ready & io_outer_release_valid;
  assign T_1942 = io_outer_release_bits_r_type == 3'h0;
  assign T_1943 = io_outer_release_bits_r_type == 3'h1;
  assign T_1944 = io_outer_release_bits_r_type == 3'h2;
  assign T_1945 = T_1942 | T_1943;
  assign T_1946 = T_1945 | T_1944;
  assign T_1947 = T_1941 & T_1946;
  assign T_1951 = T_1947 ? 8'hff : 8'h0;
  assign T_1952 = ~ T_1951;
  assign T_1954 = 8'h1 << io_outer_release_bits_addr_beat;
  assign T_1955 = ~ T_1954;
  assign T_1956 = T_1952 | T_1955;
  assign T_1957 = T_1939 & T_1956;
  assign GEN_38 = T_1922 ? T_1957 : pending_orel_data;
  assign GEN_39 = T_1646 ? 1'h1 : pending_orel_send;
  assign T_1968 = T_1946 == 1'h0;
  assign T_1970 = io_outer_release_bits_addr_beat == 3'h0;
  assign T_1971 = T_1968 | T_1970;
  assign GEN_40 = T_1971 ? 1'h1 : sending_orel;
  assign T_1983 = io_outer_release_bits_addr_beat == 3'h7;
  assign T_1984 = T_1968 | T_1983;
  assign GEN_41 = T_1984 ? 1'h0 : GEN_40;
  assign GEN_42 = T_1941 ? GEN_41 : sending_orel;
  assign GEN_43 = T_1941 ? 1'h0 : GEN_39;
  assign T_1993 = T_1941 & io_outer_release_bits_voluntary;
  assign T_2001 = T_1993 & T_1946;
  assign T_2005 = T_2003 == 3'h7;
  assign T_2007 = T_2003 + 3'h1;
  assign T_2008 = T_2007[2:0];
  assign GEN_44 = T_2001 ? T_2008 : T_2003;
  assign T_2009 = T_2001 & T_2005;
  assign T_2010 = T_1946 ? T_2003 : 3'h0;
  assign T_2011 = T_1946 ? T_2009 : T_1993;
  assign T_2012 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2014 = io_outer_grant_bits_g_type == 4'h0;
  assign T_2015 = io_outer_grant_bits_is_builtin_type & T_2014;
  assign T_2016 = T_2012 & T_2015;
  assign T_2024_0 = 3'h5;
  assign GEN_58 = {{1'd0}, T_2024_0};
  assign T_2026 = io_outer_grant_bits_g_type == GEN_58;
  assign T_2028 = io_outer_grant_bits_is_builtin_type ? T_2026 : T_2014;
  assign T_2030 = T_2016 & T_2028;
  assign T_2034 = T_2032 == 3'h7;
  assign T_2036 = T_2032 + 3'h1;
  assign T_2037 = T_2036[2:0];
  assign GEN_45 = T_2030 ? T_2037 : T_2032;
  assign T_2038 = T_2030 & T_2034;
  assign T_2039 = T_2028 ? T_2032 : 3'h0;
  assign T_2040 = T_2028 ? T_2038 : T_2016;
  assign T_2044 = T_2040 == 1'h0;
  assign T_2045 = T_2011 & T_2044;
  assign T_2047 = T_2042 + 1'h1;
  assign T_2048 = T_2047[0:0];
  assign GEN_46 = T_2045 ? T_2048 : T_2042;
  assign T_2050 = T_2011 == 1'h0;
  assign T_2051 = T_2040 & T_2050;
  assign T_2053 = T_2042 - 1'h1;
  assign T_2054 = T_2053[0:0];
  assign GEN_47 = T_2051 ? T_2054 : GEN_46;
  assign T_2056 = T_2042 > 1'h0;
  assign T_2065 = pending_orel_data >> vol_ognt_counter_up_idx;
  assign T_2066 = T_2065[0];
  assign T_2067 = T_1946 ? T_2066 : pending_orel_send;
  assign T_2068 = T_1721 & T_2067;
  assign T_2082 = T_1893_state == 2'h2;
  assign T_2083 = T_2082 ? 3'h0 : 3'h3;
  assign T_2119_addr_beat = vol_ognt_counter_up_idx;
  assign T_2119_addr_block = xact_addr_block;
  assign T_2119_client_xact_id = 2'h0;
  assign T_2119_voluntary = 1'h1;
  assign T_2119_r_type = T_2083;
  assign T_2119_data = GEN_1;
  assign GEN_1 = GEN_54;
  assign GEN_48 = 3'h1 == vol_ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_49 = 3'h2 == vol_ognt_counter_up_idx ? data_buffer_2 : GEN_48;
  assign GEN_50 = 3'h3 == vol_ognt_counter_up_idx ? data_buffer_3 : GEN_49;
  assign GEN_51 = 3'h4 == vol_ognt_counter_up_idx ? data_buffer_4 : GEN_50;
  assign GEN_52 = 3'h5 == vol_ognt_counter_up_idx ? data_buffer_5 : GEN_51;
  assign GEN_53 = 3'h6 == vol_ognt_counter_up_idx ? data_buffer_6 : GEN_52;
  assign GEN_54 = 3'h7 == vol_ognt_counter_up_idx ? data_buffer_7 : GEN_53;
  assign T_2149 = T_1656 | vol_ignt_counter_pending;
  assign T_2150 = T_2149 | scoreboard_2;
  assign T_2151 = T_2150 | vol_ognt_counter_pending;
  assign T_2153 = T_2151 == 1'h0;
  assign T_2155 = T_1721 & all_pending_done;
  assign GEN_56 = T_2155 ? 4'h0 : GEN_8;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_29 = GEN_92[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_55 = GEN_93[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_59 = GEN_94[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_60 = GEN_95[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_61 = GEN_96[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_62 = GEN_97[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_63 = GEN_98[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_64 = GEN_99[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_65 = GEN_100[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_66 = GEN_101[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_67 = GEN_102[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_68 = GEN_103[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_69 = {1{$random}};
  state = GEN_69[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_70 = {1{$random}};
  xact_addr_block = GEN_70[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_71 = {1{$random}};
  xact_vol_ir_r_type = GEN_71[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_72 = {1{$random}};
  xact_vol_ir_src = GEN_72[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_73 = {1{$random}};
  xact_vol_ir_client_xact_id = GEN_73[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_74 = {1{$random}};
  pending_irel_data = GEN_74[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_75 = {1{$random}};
  pending_orel_send = GEN_75[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_76 = {1{$random}};
  pending_orel_data = GEN_76[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_77 = {1{$random}};
  sending_orel = GEN_77[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_78 = {2{$random}};
  data_buffer_0 = GEN_78[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_79 = {2{$random}};
  data_buffer_1 = GEN_79[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_80 = {2{$random}};
  data_buffer_2 = GEN_80[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_81 = {2{$random}};
  data_buffer_3 = GEN_81[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_82 = {2{$random}};
  data_buffer_4 = GEN_82[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_83 = {2{$random}};
  data_buffer_5 = GEN_83[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_84 = {2{$random}};
  data_buffer_6 = GEN_84[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {2{$random}};
  data_buffer_7 = GEN_85[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  T_1588 = GEN_86[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_87 = {1{$random}};
  T_1619 = GEN_87[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  T_1629 = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {1{$random}};
  T_2003 = GEN_89[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {1{$random}};
  T_2032 = GEN_90[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {1{$random}};
  T_2042 = GEN_91[0:0];
  `endif
  GEN_92 = {1{$random}};
  GEN_93 = {1{$random}};
  GEN_94 = {1{$random}};
  GEN_95 = {1{$random}};
  GEN_96 = {1{$random}};
  GEN_97 = {1{$random}};
  GEN_98 = {1{$random}};
  GEN_99 = {1{$random}};
  GEN_100 = {1{$random}};
  GEN_101 = {2{$random}};
  GEN_102 = {1{$random}};
  GEN_103 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_2155) begin
        state <= 4'h0;
      end else begin
        if(T_1646) begin
          state <= 4'h7;
        end
      end
    end
    if(reset) begin
      xact_addr_block <= 26'h0;
    end else begin
      if(T_1646) begin
        xact_addr_block <= io_inner_release_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1661) begin
        if(T_1673) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_r_type <= io_inner_release_bits_r_type;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1661) begin
        if(T_1673) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_src <= io_inner_release_bits_client_id;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1661) begin
        if(T_1673) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_client_xact_id <= io_inner_release_bits_client_xact_id;
          end
        end
      end
    end
    if(reset) begin
      pending_irel_data <= 8'h0;
    end else begin
      if(T_1661) begin
        if(T_1700) begin
          pending_irel_data <= T_1717;
        end else begin
          if(T_1673) begin
            if(T_1584) begin
              pending_irel_data <= T_1696;
            end else begin
              pending_irel_data <= 8'h0;
            end
          end else begin
            if(T_1646) begin
              pending_irel_data <= 8'hff;
            end
          end
        end
      end else begin
        if(T_1646) begin
          pending_irel_data <= 8'hff;
        end
      end
    end
    if(reset) begin
      pending_orel_send <= 1'h0;
    end else begin
      if(T_1941) begin
        pending_orel_send <= 1'h0;
      end else begin
        if(T_1646) begin
          pending_orel_send <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_orel_data <= 8'h0;
    end else begin
      if(T_1922) begin
        pending_orel_data <= T_1957;
      end
    end
    if(reset) begin
      sending_orel <= 1'h0;
    end else begin
      if(T_1941) begin
        if(T_1984) begin
          sending_orel <= 1'h0;
        end else begin
          if(T_1971) begin
            sending_orel <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1544_0;
    end else begin
      if(T_1520) begin
        if(3'h0 == io_inner_release_bits_addr_beat) begin
          data_buffer_0 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1544_1;
    end else begin
      if(T_1520) begin
        if(3'h1 == io_inner_release_bits_addr_beat) begin
          data_buffer_1 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1544_2;
    end else begin
      if(T_1520) begin
        if(3'h2 == io_inner_release_bits_addr_beat) begin
          data_buffer_2 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1544_3;
    end else begin
      if(T_1520) begin
        if(3'h3 == io_inner_release_bits_addr_beat) begin
          data_buffer_3 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1544_4;
    end else begin
      if(T_1520) begin
        if(3'h4 == io_inner_release_bits_addr_beat) begin
          data_buffer_4 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1544_5;
    end else begin
      if(T_1520) begin
        if(3'h5 == io_inner_release_bits_addr_beat) begin
          data_buffer_5 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1544_6;
    end else begin
      if(T_1520) begin
        if(3'h6 == io_inner_release_bits_addr_beat) begin
          data_buffer_6 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1544_7;
    end else begin
      if(T_1520) begin
        if(3'h7 == io_inner_release_bits_addr_beat) begin
          data_buffer_7 <= GEN_0;
        end
      end
    end
    if(reset) begin
      T_1588 <= 3'h0;
    end else begin
      if(T_1586) begin
        T_1588 <= T_1593;
      end
    end
    if(reset) begin
      T_1619 <= 3'h0;
    end else begin
      if(T_1617) begin
        T_1619 <= T_1624;
      end
    end
    if(reset) begin
      T_1629 <= 1'h0;
    end else begin
      if(T_1638) begin
        T_1629 <= T_1641;
      end else begin
        if(T_1632) begin
          T_1629 <= T_1635;
        end
      end
    end
    if(reset) begin
      T_2003 <= 3'h0;
    end else begin
      if(T_2001) begin
        T_2003 <= T_2008;
      end
    end
    if(reset) begin
      T_2032 <= 3'h0;
    end else begin
      if(T_2030) begin
        T_2032 <= T_2037;
      end
    end
    if(reset) begin
      T_2042 <= 1'h0;
    end else begin
      if(T_2051) begin
        T_2042 <= T_2054;
      end else begin
        if(T_2045) begin
          T_2042 <= T_2048;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1530) begin
          $fwrite(32'h80000002,"Assertion failed: VoluntaryReleaseTracker accepted Release that wasn't voluntary!\n    at Broadcast.scala:81 assert(!(state === s_idle && io.inner.release.fire() && io.alloc.irel.should && !io.irel().isVoluntary()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1530) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_8(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_client_id,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_client_id,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [1:0] io_count
);
  reg  ram_client_xact_id [0:1];
  reg [31:0] GEN_0;
  wire  ram_client_xact_id_T_294_data;
  wire  ram_client_xact_id_T_294_addr;
  wire  ram_client_xact_id_T_294_en;
  wire  ram_client_xact_id_T_253_data;
  wire  ram_client_xact_id_T_253_addr;
  wire  ram_client_xact_id_T_253_mask;
  wire  ram_client_xact_id_T_253_en;
  reg [2:0] ram_addr_beat [0:1];
  reg [31:0] GEN_1;
  wire [2:0] ram_addr_beat_T_294_data;
  wire  ram_addr_beat_T_294_addr;
  wire  ram_addr_beat_T_294_en;
  wire [2:0] ram_addr_beat_T_253_data;
  wire  ram_addr_beat_T_253_addr;
  wire  ram_addr_beat_T_253_mask;
  wire  ram_addr_beat_T_253_en;
  reg  ram_client_id [0:1];
  reg [31:0] GEN_2;
  wire  ram_client_id_T_294_data;
  wire  ram_client_id_T_294_addr;
  wire  ram_client_id_T_294_en;
  wire  ram_client_id_T_253_data;
  wire  ram_client_id_T_253_addr;
  wire  ram_client_id_T_253_mask;
  wire  ram_client_id_T_253_en;
  reg  ram_is_builtin_type [0:1];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_294_data;
  wire  ram_is_builtin_type_T_294_addr;
  wire  ram_is_builtin_type_T_294_en;
  wire  ram_is_builtin_type_T_253_data;
  wire  ram_is_builtin_type_T_253_addr;
  wire  ram_is_builtin_type_T_253_mask;
  wire  ram_is_builtin_type_T_253_en;
  reg [2:0] ram_a_type [0:1];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_294_data;
  wire  ram_a_type_T_294_addr;
  wire  ram_a_type_T_294_en;
  wire [2:0] ram_a_type_T_253_data;
  wire  ram_a_type_T_253_addr;
  wire  ram_a_type_T_253_mask;
  wire  ram_a_type_T_253_en;
  reg  T_245;
  reg [31:0] GEN_5;
  reg  T_247;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_250;
  wire  empty;
  wire  full;
  wire  T_251;
  wire  do_enq;
  wire  T_252;
  wire  do_deq;
  wire [1:0] T_282;
  wire  T_283;
  wire  GEN_13;
  wire [1:0] T_287;
  wire  T_288;
  wire  GEN_14;
  wire  T_289;
  wire  GEN_15;
  wire  T_291;
  wire  T_293;
  wire [1:0] T_320;
  wire  ptr_diff;
  wire  T_321;
  wire [1:0] T_322;
  assign io_enq_ready = T_293;
  assign io_deq_valid = T_291;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_294_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_294_data;
  assign io_deq_bits_client_id = ram_client_id_T_294_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_294_data;
  assign io_deq_bits_a_type = ram_a_type_T_294_data;
  assign io_count = T_322;
  assign ram_client_xact_id_T_294_addr = T_247;
  assign ram_client_xact_id_T_294_en = 1'h1;
  assign ram_client_xact_id_T_294_data = ram_client_xact_id[ram_client_xact_id_T_294_addr];
  assign ram_client_xact_id_T_253_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_253_addr = T_245;
  assign ram_client_xact_id_T_253_mask = do_enq;
  assign ram_client_xact_id_T_253_en = do_enq;
  assign ram_addr_beat_T_294_addr = T_247;
  assign ram_addr_beat_T_294_en = 1'h1;
  assign ram_addr_beat_T_294_data = ram_addr_beat[ram_addr_beat_T_294_addr];
  assign ram_addr_beat_T_253_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_253_addr = T_245;
  assign ram_addr_beat_T_253_mask = do_enq;
  assign ram_addr_beat_T_253_en = do_enq;
  assign ram_client_id_T_294_addr = T_247;
  assign ram_client_id_T_294_en = 1'h1;
  assign ram_client_id_T_294_data = ram_client_id[ram_client_id_T_294_addr];
  assign ram_client_id_T_253_data = io_enq_bits_client_id;
  assign ram_client_id_T_253_addr = T_245;
  assign ram_client_id_T_253_mask = do_enq;
  assign ram_client_id_T_253_en = do_enq;
  assign ram_is_builtin_type_T_294_addr = T_247;
  assign ram_is_builtin_type_T_294_en = 1'h1;
  assign ram_is_builtin_type_T_294_data = ram_is_builtin_type[ram_is_builtin_type_T_294_addr];
  assign ram_is_builtin_type_T_253_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_253_addr = T_245;
  assign ram_is_builtin_type_T_253_mask = do_enq;
  assign ram_is_builtin_type_T_253_en = do_enq;
  assign ram_a_type_T_294_addr = T_247;
  assign ram_a_type_T_294_en = 1'h1;
  assign ram_a_type_T_294_data = ram_a_type[ram_a_type_T_294_addr];
  assign ram_a_type_T_253_data = io_enq_bits_a_type;
  assign ram_a_type_T_253_addr = T_245;
  assign ram_a_type_T_253_mask = do_enq;
  assign ram_a_type_T_253_en = do_enq;
  assign ptr_match = T_245 == T_247;
  assign T_250 = maybe_full == 1'h0;
  assign empty = ptr_match & T_250;
  assign full = ptr_match & maybe_full;
  assign T_251 = io_enq_ready & io_enq_valid;
  assign do_enq = T_251;
  assign T_252 = io_deq_ready & io_deq_valid;
  assign do_deq = T_252;
  assign T_282 = T_245 + 1'h1;
  assign T_283 = T_282[0:0];
  assign GEN_13 = do_enq ? T_283 : T_245;
  assign T_287 = T_247 + 1'h1;
  assign T_288 = T_287[0:0];
  assign GEN_14 = do_deq ? T_288 : T_247;
  assign T_289 = do_enq != do_deq;
  assign GEN_15 = T_289 ? do_enq : maybe_full;
  assign T_291 = empty == 1'h0;
  assign T_293 = full == 1'h0;
  assign T_320 = T_245 - T_247;
  assign ptr_diff = T_320[0:0];
  assign T_321 = maybe_full & ptr_match;
  assign T_322 = {T_321,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_0[0:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_1[2:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_client_id[initvar] = GEN_2[0:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  T_245 = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  T_247 = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_client_xact_id_T_253_en & ram_client_xact_id_T_253_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_253_addr] <= ram_client_xact_id_T_253_data;
    end
    if(ram_addr_beat_T_253_en & ram_addr_beat_T_253_mask) begin
      ram_addr_beat[ram_addr_beat_T_253_addr] <= ram_addr_beat_T_253_data;
    end
    if(ram_client_id_T_253_en & ram_client_id_T_253_mask) begin
      ram_client_id[ram_client_id_T_253_addr] <= ram_client_id_T_253_data;
    end
    if(ram_is_builtin_type_T_253_en & ram_is_builtin_type_T_253_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_253_addr] <= ram_is_builtin_type_T_253_data;
    end
    if(ram_a_type_T_253_en & ram_a_type_T_253_mask) begin
      ram_a_type[ram_a_type_T_253_addr] <= ram_a_type_T_253_data;
    end
    if(reset) begin
      T_245 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_245 <= T_283;
      end
    end
    if(reset) begin
      T_247 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_247 <= T_288;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_289) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module BufferedBroadcastAcquireTracker(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input   io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output  io_inner_grant_bits_client_xact_id,
  output [1:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [1:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input   io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [1:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should,
  output  io_alloc_idle,
  output [25:0] io_alloc_addr_block
);
  wire  all_pending_done;
  reg [3:0] state;
  reg [31:0] GEN_32;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_33;
  reg  xact_allocate;
  reg [31:0] GEN_41;
  reg [4:0] xact_amo_shift_bytes;
  reg [31:0] GEN_42;
  reg [4:0] xact_op_code;
  reg [31:0] GEN_43;
  reg [2:0] xact_addr_byte;
  reg [31:0] GEN_47;
  reg [1:0] xact_op_size;
  reg [31:0] GEN_78;
  wire [2:0] xact_addr_beat;
  wire  xact_iacq_client_xact_id;
  wire [2:0] xact_iacq_addr_beat;
  wire  xact_iacq_client_id;
  wire  xact_iacq_is_builtin_type;
  wire [2:0] xact_iacq_a_type;
  reg [2:0] xact_vol_ir_r_type;
  reg [31:0] GEN_79;
  reg  xact_vol_ir_src;
  reg [31:0] GEN_80;
  reg  xact_vol_ir_client_xact_id;
  reg [31:0] GEN_81;
  reg [7:0] pending_irel_data;
  reg [31:0] GEN_82;
  wire  vol_ignt_counter_pending;
  wire [2:0] vol_ignt_counter_up_idx;
  wire  vol_ignt_counter_up_done;
  wire [2:0] vol_ignt_counter_down_idx;
  wire  vol_ignt_counter_down_done;
  wire  scoreboard_6;
  wire [2:0] ignt_data_idx;
  wire  ignt_data_done;
  wire  ifin_counter_pending;
  wire [2:0] ifin_counter_up_idx;
  wire  ifin_counter_up_done;
  wire [2:0] ifin_counter_down_idx;
  wire  ifin_counter_down_done;
  reg [7:0] pending_put_data;
  reg [31:0] GEN_83;
  reg [7:0] pending_ignt_data;
  reg [31:0] GEN_84;
  wire  ognt_counter_pending;
  wire [2:0] ognt_counter_up_idx;
  wire  ognt_counter_up_done;
  wire [2:0] ognt_counter_down_idx;
  wire  ognt_counter_down_done;
  reg  pending_iprbs;
  reg [31:0] GEN_85;
  reg  pending_orel_send;
  reg [31:0] GEN_86;
  reg [7:0] pending_orel_data;
  reg [31:0] GEN_87;
  wire  vol_ognt_counter_pending;
  wire [2:0] vol_ognt_counter_up_idx;
  wire  vol_ognt_counter_up_done;
  wire [2:0] vol_ognt_counter_down_idx;
  wire  vol_ognt_counter_down_done;
  wire  T_170;
  wire  T_171;
  wire  scoreboard_3;
  reg  sending_orel;
  reg [31:0] GEN_88;
  wire  T_195_sharers;
  wire [1:0] T_241_state;
  wire  coh_inner_sharers;
  wire [1:0] coh_outer_state;
  wire  T_1611;
  wire  T_1612;
  wire  T_1613;
  wire  T_1614;
  wire [2:0] T_1623_0;
  wire  T_1625;
  wire  T_1626;
  wire  T_1627;
  wire [2:0] T_1636_0;
  wire  T_1638;
  wire  T_1639;
  wire  T_1641;
  wire  T_1643;
  wire  T_1644;
  wire  T_1646;
  wire  T_1647;
  wire  T_1649;
  wire  T_1650;
  wire  T_1652;
  wire  T_1653;
  wire  T_1654;
  wire  T_1656;
  wire  T_1658;
  wire  T_1659;
  wire  T_1660;
  wire  T_1661;
  wire  T_1663;
  wire  T_1664;
  wire  T_1666;
  wire  T_1670;
  wire  T_1671;
  wire  T_1672;
  wire  T_1674;
  wire  T_1675;
  wire  T_1677;
  wire [63:0] T_1691_0;
  wire [63:0] T_1691_1;
  wire [63:0] T_1691_2;
  wire [63:0] T_1691_3;
  wire [63:0] T_1691_4;
  wire [63:0] T_1691_5;
  wire [63:0] T_1691_6;
  wire [63:0] T_1691_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_89;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_90;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_91;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_92;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_93;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_94;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_95;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_96;
  wire [7:0] T_1709_0;
  wire [7:0] T_1709_1;
  wire [7:0] T_1709_2;
  wire [7:0] T_1709_3;
  wire [7:0] T_1709_4;
  wire [7:0] T_1709_5;
  wire [7:0] T_1709_6;
  wire [7:0] T_1709_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_97;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_98;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_99;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_100;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_101;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_102;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_103;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_104;
  wire [7:0] T_1714;
  wire  T_1716;
  wire [7:0] T_1717;
  wire  T_1719;
  wire [7:0] T_1720;
  wire  T_1722;
  wire [7:0] T_1723;
  wire  T_1725;
  wire [7:0] T_1726;
  wire  T_1728;
  wire [7:0] T_1729;
  wire  T_1731;
  wire [7:0] T_1732;
  wire  T_1734;
  wire [7:0] T_1735;
  wire  T_1737;
  wire  data_valid_0;
  wire  data_valid_1;
  wire  data_valid_2;
  wire  data_valid_3;
  wire  data_valid_4;
  wire  data_valid_5;
  wire  data_valid_6;
  wire  data_valid_7;
  wire  T_1748;
  wire  T_1749;
  wire  T_1751;
  wire  T_1752;
  wire  T_1754;
  wire  T_1755;
  wire  T_1764;
  wire  T_1765;
  wire  T_1766;
  wire  T_1767;
  wire  T_1768;
  wire  T_1769;
  wire  ignt_q_clk;
  wire  ignt_q_reset;
  wire  ignt_q_io_enq_ready;
  wire  ignt_q_io_enq_valid;
  wire  ignt_q_io_enq_bits_client_xact_id;
  wire [2:0] ignt_q_io_enq_bits_addr_beat;
  wire  ignt_q_io_enq_bits_client_id;
  wire  ignt_q_io_enq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_enq_bits_a_type;
  wire  ignt_q_io_deq_ready;
  wire  ignt_q_io_deq_valid;
  wire  ignt_q_io_deq_bits_client_xact_id;
  wire [2:0] ignt_q_io_deq_bits_addr_beat;
  wire  ignt_q_io_deq_bits_client_id;
  wire  ignt_q_io_deq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_deq_bits_a_type;
  wire [1:0] ignt_q_io_count;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [2:0] T_1812_0;
  wire  T_1814;
  wire  T_1815;
  wire  T_1817;
  wire  T_1820;
  wire  T_1821;
  wire  T_1822;
  wire  T_1823_client_xact_id;
  wire [2:0] T_1823_addr_beat;
  wire  T_1823_client_id;
  wire  T_1823_is_builtin_type;
  wire [2:0] T_1823_a_type;
  wire  T_1850;
  wire  T_1852;
  wire [2:0] T_1862_0;
  wire [2:0] T_1862_1;
  wire [2:0] T_1862_2;
  wire  T_1864;
  wire  T_1865;
  wire  T_1866;
  wire  T_1867;
  wire  T_1868;
  wire  T_1869;
  wire  T_1870;
  wire [7:0] T_1874;
  wire [7:0] T_1875;
  wire [7:0] T_1877;
  wire [7:0] T_1878;
  wire [7:0] T_1879;
  wire [7:0] T_1880;
  wire [2:0] T_1890_0;
  wire  T_1892;
  wire  T_1893;
  wire  T_1894;
  wire  T_1897;
  wire [7:0] T_1906;
  wire [7:0] T_1907;
  wire [7:0] GEN_34;
  wire [4:0] T_1915;
  wire  T_1917;
  wire  T_1918;
  wire  T_1920;
  wire  T_1921;
  wire  T_1922;
  wire [4:0] T_1923;
  wire [4:0] T_1924;
  wire [2:0] T_1925;
  wire [1:0] T_1926;
  wire [2:0] T_1939_0;
  wire [2:0] T_1939_1;
  wire [2:0] T_1939_2;
  wire  T_1941;
  wire  T_1942;
  wire  T_1943;
  wire  T_1944;
  wire  T_1945;
  wire  T_1946;
  wire  T_1947;
  wire [7:0] T_1951;
  wire [7:0] T_1952;
  wire [7:0] T_1956;
  wire [7:0] T_1958;
  wire [25:0] GEN_35;
  wire  GEN_36;
  wire [4:0] GEN_37;
  wire [4:0] GEN_38;
  wire [2:0] GEN_39;
  wire [1:0] GEN_40;
  wire [7:0] GEN_44;
  wire [7:0] GEN_45;
  wire [3:0] GEN_46;
  wire  scoreboard_0;
  wire [2:0] T_1976_0;
  wire  T_1978;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire [7:0] T_1982;
  wire  skip_outer_acquire;
  wire  T_1991;
  wire [1:0] T_1992;
  wire  T_1993;
  wire [1:0] T_1994;
  wire  T_1995;
  wire [1:0] T_1996;
  wire  T_1997;
  wire [1:0] T_1998;
  wire  T_1999;
  wire [1:0] T_2000;
  wire  T_2001;
  wire [1:0] T_2002;
  wire  T_2003;
  wire [1:0] T_2004;
  wire [1:0] T_2005;
  wire [25:0] T_2030_addr_block;
  wire [1:0] T_2030_p_type;
  wire  T_2030_client_id;
  wire  T_2055;
  wire [3:0] T_2056;
  wire  T_2065_pending;
  wire [2:0] T_2065_up_idx;
  wire  T_2065_up_done;
  wire [2:0] T_2065_down_idx;
  wire  T_2065_down_done;
  wire  T_2073;
  wire  T_2074;
  wire [1:0] T_2076;
  wire [1:0] T_2077;
  wire [1:0] GEN_410;
  wire [1:0] T_2078;
  wire [1:0] GEN_411;
  wire [1:0] T_2079;
  wire  T_2080;
  wire  T_2083;
  reg [2:0] T_2091;
  reg [31:0] GEN_105;
  wire  T_2100;
  wire  T_2103;
  wire  T_2104;
  wire  T_2105;
  wire  T_2107;
  wire  T_2108;
  wire  T_2109;
  wire  T_2110;
  wire  T_2111;
  wire  T_2113;
  reg [2:0] T_2115;
  reg [31:0] GEN_106;
  wire  T_2117;
  wire [3:0] T_2119;
  wire [2:0] T_2120;
  wire [2:0] GEN_48;
  wire  T_2121;
  wire [2:0] T_2122;
  wire  T_2123;
  reg  T_2125;
  reg [31:0] GEN_107;
  wire  T_2127;
  wire  T_2128;
  wire [1:0] T_2130;
  wire  T_2131;
  wire  GEN_49;
  wire  T_2133;
  wire  T_2134;
  wire [1:0] T_2136;
  wire  T_2137;
  wire  GEN_50;
  wire  T_2139;
  wire  T_2143;
  wire  T_2145;
  wire  T_2146;
  wire [3:0] GEN_51;
  wire  T_2150;
  wire  T_2151;
  wire  T_2156;
  wire  T_2164;
  reg [2:0] T_2166;
  reg [31:0] GEN_108;
  wire  T_2168;
  wire [3:0] T_2170;
  wire [2:0] T_2171;
  wire [2:0] GEN_52;
  wire  T_2172;
  wire [2:0] T_2173;
  wire  T_2174;
  wire  T_2175;
  wire  T_2178;
  wire  T_2179;
  wire  T_2180;
  wire  T_2181;
  wire [2:0] T_2189_0;
  wire [3:0] GEN_412;
  wire  T_2191;
  wire  T_2193;
  wire  T_2195;
  reg [2:0] T_2197;
  reg [31:0] GEN_109;
  wire  T_2199;
  wire [3:0] T_2201;
  wire [2:0] T_2202;
  wire [2:0] GEN_53;
  wire  T_2203;
  wire [2:0] T_2204;
  wire  T_2205;
  reg  T_2207;
  reg [31:0] GEN_110;
  wire  T_2209;
  wire  T_2210;
  wire [1:0] T_2212;
  wire  T_2213;
  wire  GEN_54;
  wire  T_2215;
  wire  T_2216;
  wire [1:0] T_2218;
  wire  T_2219;
  wire  GEN_55;
  wire  T_2221;
  wire  T_2223;
  wire  T_2224;
  wire [25:0] GEN_56;
  wire [7:0] GEN_57;
  wire [3:0] GEN_58;
  wire  T_2231;
  wire  T_2233;
  wire  T_2234;
  wire  T_2236;
  wire  T_2237;
  wire  T_2239;
  wire  T_2240;
  wire  T_2241;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  wire  T_2251;
  wire [7:0] T_2252;
  wire  T_2253;
  wire  T_2254;
  wire  T_2255;
  wire  T_2256;
  wire  T_2257;
  wire  T_2263;
  wire  T_2264;
  wire  T_2266;
  wire  T_2267;
  wire  T_2271;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2286;
  wire  T_2288;
  wire  T_2289;
  wire [2:0] GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  T_2303;
  wire [7:0] T_2307;
  wire [7:0] T_2308;
  wire [7:0] T_2310;
  wire [7:0] T_2311;
  wire [7:0] T_2312;
  wire [7:0] T_2314;
  wire [2:0] GEN_62;
  wire  GEN_63;
  wire  GEN_64;
  wire [7:0] GEN_65;
  wire  T_2316;
  wire [7:0] T_2333;
  wire [7:0] GEN_66;
  wire [2:0] GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire [7:0] GEN_70;
  wire  T_2334;
  wire  T_2335;
  wire  T_2337;
  wire  T_2338;
  wire  T_2339;
  wire  T_2340;
  wire  T_2341;
  wire  T_2343;
  wire  T_2344;
  wire  T_2346;
  wire  T_2347;
  wire [2:0] T_2379_addr_beat;
  wire [25:0] T_2379_addr_block;
  wire  T_2379_client_xact_id;
  wire  T_2379_voluntary;
  wire [2:0] T_2379_r_type;
  wire [63:0] T_2379_data;
  wire  T_2379_client_id;
  wire [2:0] T_2440_addr_beat;
  wire  T_2440_client_xact_id;
  wire [1:0] T_2440_manager_xact_id;
  wire  T_2440_is_builtin_type;
  wire [3:0] T_2440_g_type;
  wire [63:0] T_2440_data;
  wire  T_2440_client_id;
  wire [7:0] GEN_0;
  wire [7:0] GEN_71;
  wire [7:0] GEN_72;
  wire [7:0] GEN_73;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire  T_2521;
  wire [7:0] GEN_1;
  wire  T_2522;
  wire [7:0] GEN_2;
  wire  T_2523;
  wire [7:0] GEN_3;
  wire  T_2524;
  wire [7:0] GEN_4;
  wire  T_2525;
  wire [7:0] GEN_5;
  wire  T_2526;
  wire [7:0] GEN_6;
  wire  T_2527;
  wire [7:0] GEN_7;
  wire  T_2528;
  wire [7:0] T_2532;
  wire [7:0] T_2536;
  wire [7:0] T_2540;
  wire [7:0] T_2544;
  wire [7:0] T_2548;
  wire [7:0] T_2552;
  wire [7:0] T_2556;
  wire [7:0] T_2560;
  wire [15:0] T_2561;
  wire [15:0] T_2562;
  wire [31:0] T_2563;
  wire [15:0] T_2564;
  wire [15:0] T_2565;
  wire [31:0] T_2566;
  wire [63:0] T_2567;
  wire [63:0] T_2568;
  wire [63:0] T_2569;
  wire [63:0] GEN_8;
  wire [63:0] GEN_127;
  wire [63:0] GEN_128;
  wire [63:0] GEN_129;
  wire [63:0] GEN_130;
  wire [63:0] GEN_131;
  wire [63:0] GEN_132;
  wire [63:0] GEN_133;
  wire [63:0] T_2570;
  wire [63:0] T_2571;
  wire [63:0] GEN_9;
  wire [63:0] GEN_134;
  wire [63:0] GEN_135;
  wire [63:0] GEN_136;
  wire [63:0] GEN_137;
  wire [63:0] GEN_138;
  wire [63:0] GEN_139;
  wire [63:0] GEN_140;
  wire [63:0] GEN_141;
  wire [7:0] GEN_10;
  wire [7:0] GEN_142;
  wire [7:0] GEN_143;
  wire [7:0] GEN_144;
  wire [7:0] GEN_145;
  wire [7:0] GEN_146;
  wire [7:0] GEN_147;
  wire [7:0] GEN_148;
  wire [7:0] GEN_149;
  wire [63:0] GEN_160;
  wire [63:0] GEN_161;
  wire [63:0] GEN_162;
  wire [63:0] GEN_163;
  wire [63:0] GEN_164;
  wire [63:0] GEN_165;
  wire [63:0] GEN_166;
  wire [63:0] GEN_167;
  wire [7:0] GEN_169;
  wire [7:0] GEN_170;
  wire [7:0] GEN_171;
  wire [7:0] GEN_172;
  wire [7:0] GEN_173;
  wire [7:0] GEN_174;
  wire [7:0] GEN_175;
  wire [7:0] GEN_176;
  wire [1:0] T_2604_state;
  wire  T_2631;
  wire [7:0] T_2647;
  wire [7:0] T_2648;
  wire  T_2651;
  wire  T_2652;
  wire  T_2653;
  wire  T_2654;
  wire  T_2655;
  wire  T_2656;
  wire [7:0] T_2660;
  wire [7:0] T_2661;
  wire [7:0] T_2663;
  wire [7:0] T_2664;
  wire [7:0] T_2665;
  wire [7:0] T_2666;
  wire [7:0] GEN_177;
  wire  T_2677;
  wire  T_2679;
  wire  T_2680;
  wire  GEN_179;
  wire  T_2692;
  wire  T_2693;
  wire  GEN_180;
  wire  GEN_181;
  wire  GEN_182;
  wire  T_2702;
  wire  T_2710;
  reg [2:0] T_2712;
  reg [31:0] GEN_111;
  wire  T_2714;
  wire [3:0] T_2716;
  wire [2:0] T_2717;
  wire [2:0] GEN_183;
  wire  T_2718;
  wire [2:0] T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [2:0] T_2733_0;
  wire [3:0] GEN_413;
  wire  T_2735;
  wire  T_2737;
  wire  T_2739;
  reg [2:0] T_2741;
  reg [31:0] GEN_112;
  wire  T_2743;
  wire [3:0] T_2745;
  wire [2:0] T_2746;
  wire [2:0] GEN_184;
  wire  T_2747;
  wire [2:0] T_2748;
  wire  T_2749;
  reg  T_2751;
  reg [31:0] GEN_113;
  wire  T_2753;
  wire  T_2754;
  wire [1:0] T_2756;
  wire  T_2757;
  wire  GEN_185;
  wire  T_2759;
  wire  T_2760;
  wire [1:0] T_2762;
  wire  T_2763;
  wire  GEN_186;
  wire  T_2765;
  wire [7:0] T_2774;
  wire  T_2775;
  wire  T_2776;
  wire  T_2777;
  wire  T_2791;
  wire [2:0] T_2792;
  wire [2:0] T_2828_addr_beat;
  wire [25:0] T_2828_addr_block;
  wire [1:0] T_2828_client_xact_id;
  wire  T_2828_voluntary;
  wire [2:0] T_2828_r_type;
  wire [63:0] T_2828_data;
  wire [63:0] GEN_11;
  wire [63:0] GEN_187;
  wire [63:0] GEN_188;
  wire [63:0] GEN_189;
  wire [63:0] GEN_190;
  wire [63:0] GEN_191;
  wire [63:0] GEN_192;
  wire [63:0] GEN_193;
  wire  T_2857;
  wire  T_2860;
  wire [2:0] T_2871_0;
  wire  T_2873;
  wire  T_2874;
  wire  T_2875;
  reg [2:0] T_2877;
  reg [31:0] GEN_114;
  wire  T_2879;
  wire [3:0] T_2881;
  wire [2:0] T_2882;
  wire [2:0] GEN_195;
  wire  T_2883;
  wire [2:0] T_2884;
  wire  T_2885;
  wire  T_2891;
  wire  T_2892;
  wire [2:0] T_2900_0;
  wire [3:0] GEN_414;
  wire  T_2902;
  wire  T_2904;
  wire  T_2906;
  reg [2:0] T_2908;
  reg [31:0] GEN_115;
  wire  T_2910;
  wire [3:0] T_2912;
  wire [2:0] T_2913;
  wire [2:0] GEN_196;
  wire  T_2914;
  wire [2:0] T_2915;
  wire  T_2916;
  reg  T_2918;
  reg [31:0] GEN_116;
  wire  T_2920;
  wire  T_2921;
  wire [1:0] T_2923;
  wire  T_2924;
  wire  GEN_197;
  wire  T_2926;
  wire  T_2927;
  wire [1:0] T_2929;
  wire  T_2930;
  wire  GEN_198;
  wire  T_2932;
  wire  T_2933;
  wire [7:0] T_2937;
  wire  T_2938;
  wire  T_2940;
  wire [2:0] T_2949_0;
  wire [2:0] T_2949_1;
  wire [2:0] T_2949_2;
  wire  T_2967;
  wire  T_2968;
  wire  T_2971;
  wire  T_2972;
  wire  T_2973;
  wire  T_2974;
  wire  T_2975;
  wire  T_2976;
  wire  T_2977;
  wire  T_2978;
  wire  T_2979;
  wire  T_2980;
  wire  T_2981;
  wire [5:0] T_2984;
  wire [25:0] T_3015_addr_block;
  wire [1:0] T_3015_client_xact_id;
  wire [2:0] T_3015_addr_beat;
  wire  T_3015_is_builtin_type;
  wire [2:0] T_3015_a_type;
  wire [10:0] T_3015_union;
  wire [63:0] T_3015_data;
  wire [7:0] GEN_12;
  wire [7:0] GEN_199;
  wire [7:0] GEN_200;
  wire [7:0] GEN_201;
  wire [7:0] GEN_202;
  wire [7:0] GEN_203;
  wire [7:0] GEN_204;
  wire [7:0] GEN_205;
  wire [5:0] T_3080;
  wire [4:0] T_3081;
  wire [10:0] T_3082;
  wire [6:0] T_3084;
  wire [7:0] T_3085;
  wire [8:0] T_3087;
  wire [5:0] T_3099;
  wire [5:0] T_3101;
  wire [10:0] T_3103;
  wire [10:0] T_3105;
  wire [10:0] T_3107;
  wire [10:0] T_3109;
  wire [10:0] T_3111;
  wire [25:0] T_3140_addr_block;
  wire [1:0] T_3140_client_xact_id;
  wire [2:0] T_3140_addr_beat;
  wire  T_3140_is_builtin_type;
  wire [2:0] T_3140_a_type;
  wire [10:0] T_3140_union;
  wire [63:0] T_3140_data;
  wire [63:0] GEN_13;
  wire [63:0] GEN_206;
  wire [63:0] GEN_207;
  wire [63:0] GEN_208;
  wire [63:0] GEN_209;
  wire [63:0] GEN_210;
  wire [63:0] GEN_211;
  wire [63:0] GEN_212;
  wire [25:0] T_3168_addr_block;
  wire [1:0] T_3168_client_xact_id;
  wire [2:0] T_3168_addr_beat;
  wire  T_3168_is_builtin_type;
  wire [2:0] T_3168_a_type;
  wire [10:0] T_3168_union;
  wire [63:0] T_3168_data;
  wire  T_3197;
  wire [3:0] GEN_213;
  wire  GEN_214;
  wire [2:0] T_3207_0;
  wire [2:0] T_3207_1;
  wire [3:0] GEN_415;
  wire  T_3209;
  wire [3:0] GEN_416;
  wire  T_3210;
  wire  T_3211;
  wire  T_3213;
  wire  T_3214;
  wire [7:0] GEN_14;
  wire [7:0] GEN_215;
  wire [7:0] GEN_216;
  wire [7:0] GEN_217;
  wire [7:0] GEN_218;
  wire [7:0] GEN_219;
  wire [7:0] GEN_220;
  wire [7:0] GEN_221;
  wire  T_3215;
  wire [7:0] GEN_15;
  wire  T_3216;
  wire [7:0] GEN_16;
  wire  T_3217;
  wire [7:0] GEN_17;
  wire  T_3218;
  wire [7:0] GEN_18;
  wire  T_3219;
  wire [7:0] GEN_19;
  wire  T_3220;
  wire [7:0] GEN_20;
  wire  T_3221;
  wire [7:0] GEN_21;
  wire  T_3222;
  wire [7:0] T_3226;
  wire [7:0] T_3230;
  wire [7:0] T_3234;
  wire [7:0] T_3238;
  wire [7:0] T_3242;
  wire [7:0] T_3246;
  wire [7:0] T_3250;
  wire [7:0] T_3254;
  wire [15:0] T_3255;
  wire [15:0] T_3256;
  wire [31:0] T_3257;
  wire [15:0] T_3258;
  wire [15:0] T_3259;
  wire [31:0] T_3260;
  wire [63:0] T_3261;
  wire [63:0] T_3262;
  wire [63:0] T_3263;
  wire [63:0] GEN_22;
  wire [63:0] GEN_271;
  wire [63:0] GEN_272;
  wire [63:0] GEN_273;
  wire [63:0] GEN_274;
  wire [63:0] GEN_275;
  wire [63:0] GEN_276;
  wire [63:0] GEN_277;
  wire [63:0] T_3264;
  wire [63:0] T_3265;
  wire [63:0] GEN_23;
  wire [63:0] GEN_278;
  wire [63:0] GEN_279;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [7:0] GEN_24;
  wire [7:0] GEN_286;
  wire [7:0] GEN_287;
  wire [7:0] GEN_288;
  wire [7:0] GEN_289;
  wire [7:0] GEN_290;
  wire [7:0] GEN_291;
  wire [7:0] GEN_292;
  wire [7:0] GEN_293;
  wire [63:0] GEN_304;
  wire [63:0] GEN_305;
  wire [63:0] GEN_306;
  wire [63:0] GEN_307;
  wire [63:0] GEN_308;
  wire [63:0] GEN_309;
  wire [63:0] GEN_310;
  wire [63:0] GEN_311;
  wire [7:0] GEN_313;
  wire [7:0] GEN_314;
  wire [7:0] GEN_315;
  wire [7:0] GEN_316;
  wire [7:0] GEN_317;
  wire [7:0] GEN_318;
  wire [7:0] GEN_319;
  wire [7:0] GEN_320;
  wire  T_3268;
  wire  T_3269;
  wire  T_3281;
  wire  T_3283;
  wire [2:0] T_3291_0;
  wire [3:0] GEN_417;
  wire  T_3293;
  wire  T_3295;
  wire  T_3297;
  reg [2:0] T_3299;
  reg [31:0] GEN_117;
  wire  T_3301;
  wire [3:0] T_3303;
  wire [2:0] T_3304;
  wire [2:0] GEN_321;
  wire  T_3305;
  wire [2:0] T_3306;
  wire  T_3307;
  wire  T_3308;
  reg [2:0] T_3314;
  reg [31:0] GEN_118;
  reg  T_3324;
  reg [31:0] GEN_119;
  wire  T_3326;
  wire  T_3327;
  wire [1:0] T_3329;
  wire  T_3330;
  wire  GEN_323;
  wire  T_3332;
  wire  T_3333;
  wire [1:0] T_3335;
  wire  T_3336;
  wire  GEN_324;
  wire  T_3338;
  wire  T_3343;
  wire [7:0] T_3360;
  wire [2:0] T_3370_0;
  wire [2:0] T_3370_1;
  wire [3:0] GEN_418;
  wire  T_3372;
  wire [3:0] GEN_419;
  wire  T_3373;
  wire  T_3374;
  wire  T_3376;
  wire  T_3377;
  wire [7:0] T_3382;
  wire [7:0] T_3384;
  wire [7:0] T_3385;
  wire [7:0] T_3386;
  wire [7:0] GEN_327;
  wire  T_3389;
  wire  T_3390;
  wire  T_3393;
  wire  T_3395;
  wire  T_3412;
  wire [2:0] T_3413;
  wire  T_3414;
  wire [2:0] T_3415;
  wire  T_3416;
  wire [2:0] T_3417;
  wire  T_3418;
  wire [2:0] T_3419;
  wire  T_3420;
  wire [2:0] T_3421;
  wire  T_3422;
  wire [2:0] T_3423;
  wire  T_3424;
  wire [2:0] T_3425;
  wire [2:0] T_3426;
  wire [2:0] T_3455_addr_beat;
  wire  T_3455_client_xact_id;
  wire [1:0] T_3455_manager_xact_id;
  wire  T_3455_is_builtin_type;
  wire [3:0] T_3455_g_type;
  wire [63:0] T_3455_data;
  wire  T_3455_client_id;
  wire [63:0] GEN_25;
  wire [63:0] GEN_328;
  wire [63:0] GEN_329;
  wire [63:0] GEN_330;
  wire [63:0] GEN_331;
  wire [63:0] GEN_332;
  wire [63:0] GEN_333;
  wire [63:0] GEN_334;
  wire [2:0] T_3491_0;
  wire [3:0] GEN_420;
  wire  T_3493;
  wire  T_3495;
  wire  T_3497;
  reg [2:0] T_3499;
  reg [31:0] GEN_120;
  wire  T_3501;
  wire [3:0] T_3503;
  wire [2:0] T_3504;
  wire [2:0] GEN_335;
  wire  T_3505;
  wire [2:0] T_3506;
  wire  T_3507;
  wire  T_3512;
  wire  T_3514;
  wire [2:0] T_3522_0;
  wire [2:0] T_3522_1;
  wire [3:0] GEN_421;
  wire  T_3524;
  wire [3:0] GEN_422;
  wire  T_3525;
  wire  T_3526;
  wire  T_3528;
  wire [7:0] T_3529;
  wire  T_3530;
  wire  T_3532;
  wire  T_3533;
  wire  GEN_338;
  wire  GEN_339;
  wire [2:0] GEN_340;
  wire  GEN_341;
  wire [1:0] GEN_342;
  wire  GEN_343;
  wire [3:0] GEN_344;
  wire [63:0] GEN_345;
  wire  GEN_346;
  wire  GEN_349;
  wire  T_3540;
  wire [1:0] GEN_350;
  wire  T_3551;
  wire  T_3552;
  wire [2:0] T_3562_0;
  wire [2:0] T_3562_1;
  wire [2:0] T_3562_2;
  wire  T_3564;
  wire  T_3565;
  wire  T_3566;
  wire  T_3567;
  wire  T_3568;
  wire  T_3569;
  wire  T_3570;
  wire  T_3571;
  wire  T_3573;
  wire  T_3574;
  wire  T_3603;
  wire [7:0] T_3604;
  wire [7:0] T_3606;
  wire [7:0] T_3607;
  wire  T_3608;
  wire  T_3609;
  wire  T_3610;
  wire  T_3611;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3615;
  wire [7:0] T_3619;
  wire [7:0] T_3623;
  wire [7:0] T_3627;
  wire [7:0] T_3631;
  wire [7:0] T_3635;
  wire [7:0] T_3639;
  wire [7:0] T_3643;
  wire [7:0] T_3647;
  wire [15:0] T_3648;
  wire [15:0] T_3649;
  wire [31:0] T_3650;
  wire [15:0] T_3651;
  wire [15:0] T_3652;
  wire [31:0] T_3653;
  wire [63:0] T_3654;
  wire [63:0] T_3655;
  wire [63:0] GEN_26;
  wire [63:0] GEN_351;
  wire [63:0] GEN_352;
  wire [63:0] GEN_353;
  wire [63:0] GEN_354;
  wire [63:0] GEN_355;
  wire [63:0] GEN_356;
  wire [63:0] GEN_357;
  wire [63:0] T_3656;
  wire [63:0] T_3657;
  wire [63:0] T_3658;
  wire [63:0] GEN_27;
  wire [63:0] GEN_358;
  wire [63:0] GEN_359;
  wire [63:0] GEN_360;
  wire [63:0] GEN_361;
  wire [63:0] GEN_362;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [7:0] GEN_28;
  wire [7:0] GEN_366;
  wire [7:0] GEN_367;
  wire [7:0] GEN_368;
  wire [7:0] GEN_369;
  wire [7:0] GEN_370;
  wire [7:0] GEN_371;
  wire [7:0] GEN_372;
  wire [7:0] T_3695;
  wire [7:0] GEN_29;
  wire [7:0] GEN_373;
  wire [7:0] GEN_374;
  wire [7:0] GEN_375;
  wire [7:0] GEN_376;
  wire [7:0] GEN_377;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [63:0] GEN_383;
  wire [63:0] GEN_384;
  wire [63:0] GEN_385;
  wire [63:0] GEN_386;
  wire [63:0] GEN_387;
  wire [63:0] GEN_388;
  wire [63:0] GEN_389;
  wire [63:0] GEN_390;
  wire [7:0] GEN_393;
  wire [7:0] GEN_394;
  wire [7:0] GEN_395;
  wire [7:0] GEN_396;
  wire [7:0] GEN_397;
  wire [7:0] GEN_398;
  wire [7:0] GEN_399;
  wire [7:0] GEN_400;
  wire  T_3698;
  wire  T_3699;
  wire  T_3700;
  wire  T_3701;
  wire  T_3702;
  wire  T_3703;
  wire  T_3704;
  wire  T_3706;
  wire  T_3708;
  wire [3:0] GEN_401;
  wire [7:0] GEN_402;
  wire [7:0] GEN_403;
  wire [7:0] GEN_404;
  wire [7:0] GEN_405;
  wire [7:0] GEN_406;
  wire [7:0] GEN_407;
  wire [7:0] GEN_408;
  wire [7:0] GEN_409;
  wire  GEN_30;
  reg [31:0] GEN_121;
  wire  GEN_31;
  reg [31:0] GEN_122;
  Queue_8 ignt_q (
    .clk(ignt_q_clk),
    .reset(ignt_q_reset),
    .io_enq_ready(ignt_q_io_enq_ready),
    .io_enq_valid(ignt_q_io_enq_valid),
    .io_enq_bits_client_xact_id(ignt_q_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(ignt_q_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(ignt_q_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(ignt_q_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(ignt_q_io_enq_bits_a_type),
    .io_deq_ready(ignt_q_io_deq_ready),
    .io_deq_valid(ignt_q_io_deq_valid),
    .io_deq_bits_client_xact_id(ignt_q_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(ignt_q_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(ignt_q_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(ignt_q_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(ignt_q_io_deq_bits_a_type),
    .io_count(ignt_q_io_count)
  );
  assign io_inner_acquire_ready = T_1981;
  assign io_inner_grant_valid = GEN_349;
  assign io_inner_grant_bits_addr_beat = GEN_340;
  assign io_inner_grant_bits_client_xact_id = GEN_341;
  assign io_inner_grant_bits_manager_xact_id = GEN_342;
  assign io_inner_grant_bits_is_builtin_type = GEN_343;
  assign io_inner_grant_bits_g_type = GEN_344;
  assign io_inner_grant_bits_data = GEN_345;
  assign io_inner_grant_bits_client_id = GEN_346;
  assign io_inner_finish_ready = T_2337;
  assign io_inner_probe_valid = T_2083;
  assign io_inner_probe_bits_addr_block = T_2030_addr_block;
  assign io_inner_probe_bits_p_type = T_2030_p_type;
  assign io_inner_probe_bits_client_id = T_2030_client_id;
  assign io_inner_release_ready = T_2274;
  assign io_outer_acquire_valid = T_2968;
  assign io_outer_acquire_bits_addr_block = T_3168_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3168_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3168_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3168_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3168_a_type;
  assign io_outer_acquire_bits_union = T_3168_union;
  assign io_outer_acquire_bits_data = T_3168_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2777;
  assign io_outer_release_bits_addr_beat = T_2828_addr_beat;
  assign io_outer_release_bits_addr_block = T_2828_addr_block;
  assign io_outer_release_bits_client_xact_id = T_2828_client_xact_id;
  assign io_outer_release_bits_voluntary = T_2828_voluntary;
  assign io_outer_release_bits_r_type = T_2828_r_type;
  assign io_outer_release_bits_data = T_2828_data;
  assign io_outer_grant_ready = GEN_214;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_30;
  assign io_outer_finish_bits_manager_id = GEN_31;
  assign io_alloc_iacq_matches = T_1749;
  assign io_alloc_iacq_can = T_1611;
  assign io_alloc_irel_matches = T_1752;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1755;
  assign io_alloc_oprb_can = 1'h0;
  assign io_alloc_idle = T_1611;
  assign io_alloc_addr_block = xact_addr_block;
  assign all_pending_done = T_3706;
  assign xact_addr_beat = xact_iacq_addr_beat;
  assign xact_iacq_client_xact_id = T_1823_client_xact_id;
  assign xact_iacq_addr_beat = T_1823_addr_beat;
  assign xact_iacq_client_id = T_1823_client_id;
  assign xact_iacq_is_builtin_type = T_1823_is_builtin_type;
  assign xact_iacq_a_type = T_1823_a_type;
  assign vol_ignt_counter_pending = T_2221;
  assign vol_ignt_counter_up_idx = T_2173;
  assign vol_ignt_counter_up_done = T_2174;
  assign vol_ignt_counter_down_idx = T_2204;
  assign vol_ignt_counter_down_done = T_2205;
  assign scoreboard_6 = T_1850;
  assign ignt_data_idx = T_3506;
  assign ignt_data_done = T_3507;
  assign ifin_counter_pending = T_3338;
  assign ifin_counter_up_idx = T_3306;
  assign ifin_counter_up_done = T_3307;
  assign ifin_counter_down_idx = 3'h0;
  assign ifin_counter_down_done = T_3308;
  assign ognt_counter_pending = T_2932;
  assign ognt_counter_up_idx = T_2884;
  assign ognt_counter_up_done = T_2885;
  assign ognt_counter_down_idx = T_2915;
  assign ognt_counter_down_done = T_2916;
  assign vol_ognt_counter_pending = T_2765;
  assign vol_ognt_counter_up_idx = T_2719;
  assign vol_ognt_counter_up_done = T_2720;
  assign vol_ognt_counter_down_idx = T_2748;
  assign vol_ognt_counter_down_done = T_2749;
  assign T_170 = pending_orel_data != 8'h0;
  assign T_171 = pending_orel_send | T_170;
  assign scoreboard_3 = T_171 | vol_ognt_counter_pending;
  assign T_195_sharers = 1'h0;
  assign T_241_state = 2'h0;
  assign coh_inner_sharers = T_195_sharers;
  assign coh_outer_state = T_241_state;
  assign T_1611 = state == 4'h0;
  assign T_1612 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1613 = T_1611 & T_1612;
  assign T_1614 = T_1613 & io_alloc_iacq_should;
  assign T_1623_0 = 3'h3;
  assign T_1625 = io_inner_acquire_bits_a_type == T_1623_0;
  assign T_1626 = io_inner_acquire_bits_is_builtin_type & T_1625;
  assign T_1627 = T_1614 & T_1626;
  assign T_1636_0 = 3'h3;
  assign T_1638 = io_inner_acquire_bits_a_type == T_1636_0;
  assign T_1639 = io_inner_acquire_bits_is_builtin_type & T_1638;
  assign T_1641 = T_1639 == 1'h0;
  assign T_1643 = io_inner_acquire_bits_addr_beat == 3'h0;
  assign T_1644 = T_1641 | T_1643;
  assign T_1646 = T_1644 == 1'h0;
  assign T_1647 = T_1627 & T_1646;
  assign T_1649 = T_1647 == 1'h0;
  assign T_1650 = T_1649 | reset;
  assign T_1652 = T_1650 == 1'h0;
  assign T_1653 = state != 4'h0;
  assign T_1654 = T_1653 & scoreboard_6;
  assign T_1656 = xact_iacq_a_type == 3'h5;
  assign T_1658 = xact_iacq_a_type == 3'h6;
  assign T_1659 = T_1656 | T_1658;
  assign T_1660 = xact_iacq_is_builtin_type & T_1659;
  assign T_1661 = T_1654 & T_1660;
  assign T_1663 = T_1661 == 1'h0;
  assign T_1664 = T_1663 | reset;
  assign T_1666 = T_1664 == 1'h0;
  assign T_1670 = xact_iacq_a_type == 3'h4;
  assign T_1671 = xact_iacq_is_builtin_type & T_1670;
  assign T_1672 = T_1654 & T_1671;
  assign T_1674 = T_1672 == 1'h0;
  assign T_1675 = T_1674 | reset;
  assign T_1677 = T_1675 == 1'h0;
  assign T_1691_0 = 64'h0;
  assign T_1691_1 = 64'h0;
  assign T_1691_2 = 64'h0;
  assign T_1691_3 = 64'h0;
  assign T_1691_4 = 64'h0;
  assign T_1691_5 = 64'h0;
  assign T_1691_6 = 64'h0;
  assign T_1691_7 = 64'h0;
  assign T_1709_0 = 8'h0;
  assign T_1709_1 = 8'h0;
  assign T_1709_2 = 8'h0;
  assign T_1709_3 = 8'h0;
  assign T_1709_4 = 8'h0;
  assign T_1709_5 = 8'h0;
  assign T_1709_6 = 8'h0;
  assign T_1709_7 = 8'h0;
  assign T_1714 = ~ wmask_buffer_0;
  assign T_1716 = T_1714 == 8'h0;
  assign T_1717 = ~ wmask_buffer_1;
  assign T_1719 = T_1717 == 8'h0;
  assign T_1720 = ~ wmask_buffer_2;
  assign T_1722 = T_1720 == 8'h0;
  assign T_1723 = ~ wmask_buffer_3;
  assign T_1725 = T_1723 == 8'h0;
  assign T_1726 = ~ wmask_buffer_4;
  assign T_1728 = T_1726 == 8'h0;
  assign T_1729 = ~ wmask_buffer_5;
  assign T_1731 = T_1729 == 8'h0;
  assign T_1732 = ~ wmask_buffer_6;
  assign T_1734 = T_1732 == 8'h0;
  assign T_1735 = ~ wmask_buffer_7;
  assign T_1737 = T_1735 == 8'h0;
  assign data_valid_0 = T_1716;
  assign data_valid_1 = T_1719;
  assign data_valid_2 = T_1722;
  assign data_valid_3 = T_1725;
  assign data_valid_4 = T_1728;
  assign data_valid_5 = T_1731;
  assign data_valid_6 = T_1734;
  assign data_valid_7 = T_1737;
  assign T_1748 = io_inner_acquire_bits_addr_block == xact_addr_block;
  assign T_1749 = T_1653 & T_1748;
  assign T_1751 = io_inner_release_bits_addr_block == xact_addr_block;
  assign T_1752 = T_1653 & T_1751;
  assign T_1754 = io_outer_probe_bits_addr_block == xact_addr_block;
  assign T_1755 = T_1653 & T_1754;
  assign T_1764 = xact_iacq_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1765 = xact_iacq_client_id == io_inner_acquire_bits_client_id;
  assign T_1766 = T_1764 & T_1765;
  assign T_1767 = T_1766 & scoreboard_6;
  assign T_1768 = xact_iacq_addr_beat == io_inner_acquire_bits_addr_beat;
  assign T_1769 = T_1767 & T_1768;
  assign ignt_q_clk = clk;
  assign ignt_q_reset = reset;
  assign ignt_q_io_enq_valid = T_1822;
  assign ignt_q_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign ignt_q_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign ignt_q_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign ignt_q_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign ignt_q_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign ignt_q_io_deq_ready = GEN_339;
  assign T_1797 = T_1611 & io_alloc_iacq_should;
  assign T_1798 = T_1797 & io_inner_acquire_valid;
  assign T_1800 = T_1769 == 1'h0;
  assign T_1801 = T_1800 & scoreboard_6;
  assign T_1803 = T_1801 & T_1612;
  assign T_1812_0 = 3'h3;
  assign T_1814 = io_inner_acquire_bits_a_type == T_1812_0;
  assign T_1815 = io_inner_acquire_bits_is_builtin_type & T_1814;
  assign T_1817 = T_1815 == 1'h0;
  assign T_1820 = T_1817 | T_1643;
  assign T_1821 = T_1803 & T_1820;
  assign T_1822 = T_1798 | T_1821;
  assign T_1823_client_xact_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_xact_id : ignt_q_io_enq_bits_client_xact_id;
  assign T_1823_addr_beat = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_addr_beat : ignt_q_io_enq_bits_addr_beat;
  assign T_1823_client_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_id : ignt_q_io_enq_bits_client_id;
  assign T_1823_is_builtin_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_is_builtin_type : ignt_q_io_enq_bits_is_builtin_type;
  assign T_1823_a_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_a_type : ignt_q_io_enq_bits_a_type;
  assign T_1850 = ignt_q_io_count > 2'h0;
  assign T_1852 = T_1653 | io_alloc_iacq_should;
  assign T_1862_0 = 3'h2;
  assign T_1862_1 = 3'h3;
  assign T_1862_2 = 3'h4;
  assign T_1864 = io_inner_acquire_bits_a_type == T_1862_0;
  assign T_1865 = io_inner_acquire_bits_a_type == T_1862_1;
  assign T_1866 = io_inner_acquire_bits_a_type == T_1862_2;
  assign T_1867 = T_1864 | T_1865;
  assign T_1868 = T_1867 | T_1866;
  assign T_1869 = io_inner_acquire_bits_is_builtin_type & T_1868;
  assign T_1870 = T_1612 & T_1869;
  assign T_1874 = T_1870 ? 8'hff : 8'h0;
  assign T_1875 = ~ T_1874;
  assign T_1877 = 8'h1 << io_inner_acquire_bits_addr_beat;
  assign T_1878 = ~ T_1877;
  assign T_1879 = T_1875 | T_1878;
  assign T_1880 = pending_put_data & T_1879;
  assign T_1890_0 = 3'h3;
  assign T_1892 = io_inner_acquire_bits_a_type == T_1890_0;
  assign T_1893 = io_inner_acquire_bits_is_builtin_type & T_1892;
  assign T_1894 = T_1612 & T_1893;
  assign T_1897 = T_1894 & T_1643;
  assign T_1906 = T_1897 ? 8'hfe : 8'h0;
  assign T_1907 = T_1880 | T_1906;
  assign GEN_34 = T_1852 ? T_1907 : pending_put_data;
  assign T_1915 = 4'h8 * 4'h0;
  assign T_1917 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1918 = io_inner_acquire_bits_is_builtin_type & T_1917;
  assign T_1920 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1921 = io_inner_acquire_bits_is_builtin_type & T_1920;
  assign T_1922 = T_1918 | T_1921;
  assign T_1923 = io_inner_acquire_bits_union[5:1];
  assign T_1924 = T_1922 ? 5'h1 : T_1923;
  assign T_1925 = io_inner_acquire_bits_union[10:8];
  assign T_1926 = io_inner_acquire_bits_union[7:6];
  assign T_1939_0 = 3'h2;
  assign T_1939_1 = 3'h3;
  assign T_1939_2 = 3'h4;
  assign T_1941 = io_inner_acquire_bits_a_type == T_1939_0;
  assign T_1942 = io_inner_acquire_bits_a_type == T_1939_1;
  assign T_1943 = io_inner_acquire_bits_a_type == T_1939_2;
  assign T_1944 = T_1941 | T_1942;
  assign T_1945 = T_1944 | T_1943;
  assign T_1946 = io_inner_acquire_bits_is_builtin_type & T_1945;
  assign T_1947 = T_1612 & T_1946;
  assign T_1951 = T_1947 ? 8'hff : 8'h0;
  assign T_1952 = ~ T_1951;
  assign T_1956 = T_1952 | T_1878;
  assign T_1958 = T_1921 ? T_1956 : 8'h0;
  assign GEN_35 = T_1798 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_36 = T_1798 ? 1'h0 : xact_allocate;
  assign GEN_37 = T_1798 ? T_1915 : xact_amo_shift_bytes;
  assign GEN_38 = T_1798 ? T_1924 : xact_op_code;
  assign GEN_39 = T_1798 ? T_1925 : xact_addr_byte;
  assign GEN_40 = T_1798 ? T_1926 : xact_op_size;
  assign GEN_44 = T_1798 ? T_1958 : GEN_34;
  assign GEN_45 = T_1798 ? 8'h0 : pending_ignt_data;
  assign GEN_46 = T_1798 ? 4'h5 : state;
  assign scoreboard_0 = pending_put_data != 8'h0;
  assign T_1976_0 = 3'h3;
  assign T_1978 = io_inner_acquire_bits_a_type == T_1976_0;
  assign T_1979 = io_inner_acquire_bits_is_builtin_type & T_1978;
  assign T_1980 = T_1767 & T_1979;
  assign T_1981 = T_1611 | T_1980;
  assign T_1982 = ~ pending_ignt_data;
  assign skip_outer_acquire = T_1982 == 8'h0;
  assign T_1991 = 3'h4 == xact_iacq_a_type;
  assign T_1992 = T_1991 ? 2'h0 : 2'h2;
  assign T_1993 = 3'h6 == xact_iacq_a_type;
  assign T_1994 = T_1993 ? 2'h0 : T_1992;
  assign T_1995 = 3'h5 == xact_iacq_a_type;
  assign T_1996 = T_1995 ? 2'h2 : T_1994;
  assign T_1997 = 3'h2 == xact_iacq_a_type;
  assign T_1998 = T_1997 ? 2'h0 : T_1996;
  assign T_1999 = 3'h0 == xact_iacq_a_type;
  assign T_2000 = T_1999 ? 2'h2 : T_1998;
  assign T_2001 = 3'h3 == xact_iacq_a_type;
  assign T_2002 = T_2001 ? 2'h0 : T_2000;
  assign T_2003 = 3'h1 == xact_iacq_a_type;
  assign T_2004 = T_2003 ? 2'h2 : T_2002;
  assign T_2005 = xact_iacq_is_builtin_type ? T_2004 : 2'h0;
  assign T_2030_addr_block = xact_addr_block;
  assign T_2030_p_type = T_2005;
  assign T_2030_client_id = 1'h0;
  assign T_2055 = skip_outer_acquire == 1'h0;
  assign T_2056 = T_2055 ? 4'h6 : 4'h7;
  assign T_2065_pending = T_2139;
  assign T_2065_up_idx = 3'h0;
  assign T_2065_up_done = T_2073;
  assign T_2065_down_idx = T_2122;
  assign T_2065_down_done = T_2123;
  assign T_2073 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2074 = ~ T_2073;
  assign T_2076 = 2'h1 << io_inner_probe_bits_client_id;
  assign T_2077 = ~ T_2076;
  assign GEN_410 = {{1'd0}, T_2074};
  assign T_2078 = GEN_410 | T_2077;
  assign GEN_411 = {{1'd0}, pending_iprbs};
  assign T_2079 = GEN_411 & T_2078;
  assign T_2080 = state == 4'h5;
  assign T_2083 = T_2080 & pending_iprbs;
  assign T_2100 = io_inner_release_ready & io_inner_release_valid;
  assign T_2103 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2104 = T_1653 & T_2103;
  assign T_2105 = T_2100 & T_2104;
  assign T_2107 = io_inner_release_bits_r_type == 3'h0;
  assign T_2108 = io_inner_release_bits_r_type == 3'h1;
  assign T_2109 = io_inner_release_bits_r_type == 3'h2;
  assign T_2110 = T_2107 | T_2108;
  assign T_2111 = T_2110 | T_2109;
  assign T_2113 = T_2105 & T_2111;
  assign T_2117 = T_2115 == 3'h7;
  assign T_2119 = T_2115 + 3'h1;
  assign T_2120 = T_2119[2:0];
  assign GEN_48 = T_2113 ? T_2120 : T_2115;
  assign T_2121 = T_2113 & T_2117;
  assign T_2122 = T_2111 ? T_2115 : 3'h0;
  assign T_2123 = T_2111 ? T_2121 : T_2105;
  assign T_2127 = T_2123 == 1'h0;
  assign T_2128 = T_2073 & T_2127;
  assign T_2130 = T_2125 + 1'h1;
  assign T_2131 = T_2130[0:0];
  assign GEN_49 = T_2128 ? T_2131 : T_2125;
  assign T_2133 = T_2073 == 1'h0;
  assign T_2134 = T_2123 & T_2133;
  assign T_2136 = T_2125 - 1'h1;
  assign T_2137 = T_2136[0:0];
  assign GEN_50 = T_2134 ? T_2137 : GEN_49;
  assign T_2139 = T_2125 > 1'h0;
  assign T_2143 = pending_iprbs | T_2065_pending;
  assign T_2145 = T_2143 == 1'h0;
  assign T_2146 = T_2080 & T_2145;
  assign GEN_51 = T_2146 ? T_2056 : GEN_46;
  assign T_2150 = T_1611 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2151 = T_2150 & io_inner_release_bits_voluntary;
  assign T_2156 = T_2100 & T_2151;
  assign T_2164 = T_2156 & T_2111;
  assign T_2168 = T_2166 == 3'h7;
  assign T_2170 = T_2166 + 3'h1;
  assign T_2171 = T_2170[2:0];
  assign GEN_52 = T_2164 ? T_2171 : T_2166;
  assign T_2172 = T_2164 & T_2168;
  assign T_2173 = T_2111 ? T_2166 : 3'h0;
  assign T_2174 = T_2111 ? T_2172 : T_2156;
  assign T_2175 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_2178 = io_inner_grant_bits_g_type == 4'h0;
  assign T_2179 = io_inner_grant_bits_is_builtin_type & T_2178;
  assign T_2180 = T_1653 & T_2179;
  assign T_2181 = T_2175 & T_2180;
  assign T_2189_0 = 3'h5;
  assign GEN_412 = {{1'd0}, T_2189_0};
  assign T_2191 = io_inner_grant_bits_g_type == GEN_412;
  assign T_2193 = io_inner_grant_bits_is_builtin_type ? T_2191 : T_2178;
  assign T_2195 = T_2181 & T_2193;
  assign T_2199 = T_2197 == 3'h7;
  assign T_2201 = T_2197 + 3'h1;
  assign T_2202 = T_2201[2:0];
  assign GEN_53 = T_2195 ? T_2202 : T_2197;
  assign T_2203 = T_2195 & T_2199;
  assign T_2204 = T_2193 ? T_2197 : 3'h0;
  assign T_2205 = T_2193 ? T_2203 : T_2181;
  assign T_2209 = T_2205 == 1'h0;
  assign T_2210 = T_2174 & T_2209;
  assign T_2212 = T_2207 + 1'h1;
  assign T_2213 = T_2212[0:0];
  assign GEN_54 = T_2210 ? T_2213 : T_2207;
  assign T_2215 = T_2174 == 1'h0;
  assign T_2216 = T_2205 & T_2215;
  assign T_2218 = T_2207 - 1'h1;
  assign T_2219 = T_2218[0:0];
  assign GEN_55 = T_2216 ? T_2219 : GEN_54;
  assign T_2221 = T_2207 > 1'h0;
  assign T_2223 = T_1611 & io_alloc_irel_should;
  assign T_2224 = T_2223 & io_inner_release_valid;
  assign GEN_56 = T_2224 ? io_inner_release_bits_addr_block : GEN_35;
  assign GEN_57 = T_2224 ? 8'hff : pending_irel_data;
  assign GEN_58 = T_2224 ? 4'h7 : GEN_51;
  assign T_2231 = T_1751 & io_inner_release_bits_voluntary;
  assign T_2233 = state == 4'h8;
  assign T_2234 = T_1611 | T_2233;
  assign T_2236 = T_2234 == 1'h0;
  assign T_2237 = T_2231 & T_2236;
  assign T_2239 = all_pending_done == 1'h0;
  assign T_2240 = T_2237 & T_2239;
  assign T_2241 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2243 = T_2241 == 1'h0;
  assign T_2244 = T_2240 & T_2243;
  assign T_2247 = T_2175 == 1'h0;
  assign T_2248 = T_2244 & T_2247;
  assign T_2250 = vol_ignt_counter_pending == 1'h0;
  assign T_2251 = T_2248 & T_2250;
  assign T_2252 = pending_orel_data >> io_inner_release_bits_addr_beat;
  assign T_2253 = T_2252[0];
  assign T_2254 = sending_orel & T_2253;
  assign T_2255 = io_outer_release_ready & io_outer_release_valid;
  assign T_2256 = io_inner_release_bits_addr_beat == io_outer_release_bits_addr_beat;
  assign T_2257 = T_2255 & T_2256;
  assign T_2263 = T_2254 | T_2257;
  assign T_2264 = T_2111 & T_2263;
  assign T_2266 = T_2264 == 1'h0;
  assign T_2267 = T_2251 & T_2266;
  assign T_2271 = T_1751 & T_2103;
  assign T_2273 = T_2271 & T_2080;
  assign T_2274 = T_2267 | T_2273;
  assign T_2275 = T_2274 & io_inner_release_valid;
  assign T_2276 = T_2224 | T_2275;
  assign T_2277 = T_2276 & io_inner_release_ready;
  assign T_2286 = T_2111 == 1'h0;
  assign T_2288 = io_inner_release_bits_addr_beat == 3'h0;
  assign T_2289 = T_2286 | T_2288;
  assign GEN_59 = io_inner_release_bits_voluntary ? io_inner_release_bits_r_type : xact_vol_ir_r_type;
  assign GEN_60 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_id : xact_vol_ir_src;
  assign GEN_61 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_xact_id : xact_vol_ir_client_xact_id;
  assign T_2303 = T_2100 & T_2111;
  assign T_2307 = T_2303 ? 8'hff : 8'h0;
  assign T_2308 = ~ T_2307;
  assign T_2310 = 8'h1 << io_inner_release_bits_addr_beat;
  assign T_2311 = ~ T_2310;
  assign T_2312 = T_2308 | T_2311;
  assign T_2314 = T_2111 ? T_2312 : 8'h0;
  assign GEN_62 = T_2289 ? GEN_59 : xact_vol_ir_r_type;
  assign GEN_63 = T_2289 ? GEN_60 : xact_vol_ir_src;
  assign GEN_64 = T_2289 ? GEN_61 : xact_vol_ir_client_xact_id;
  assign GEN_65 = T_2289 ? T_2314 : GEN_57;
  assign T_2316 = T_2289 == 1'h0;
  assign T_2333 = pending_irel_data & T_2312;
  assign GEN_66 = T_2316 ? T_2333 : GEN_65;
  assign GEN_67 = T_2277 ? GEN_62 : xact_vol_ir_r_type;
  assign GEN_68 = T_2277 ? GEN_63 : xact_vol_ir_src;
  assign GEN_69 = T_2277 ? GEN_64 : xact_vol_ir_client_xact_id;
  assign GEN_70 = T_2277 ? GEN_66 : GEN_57;
  assign T_2334 = state == 4'h3;
  assign T_2335 = state == 4'h4;
  assign T_2337 = state == 4'h7;
  assign T_2338 = T_2334 | T_2335;
  assign T_2339 = T_2338 | T_2080;
  assign T_2340 = T_2339 | T_2337;
  assign T_2341 = T_2340 & vol_ignt_counter_pending;
  assign T_2343 = pending_irel_data != 8'h0;
  assign T_2344 = T_2343 | vol_ognt_counter_pending;
  assign T_2346 = T_2344 == 1'h0;
  assign T_2347 = T_2341 & T_2346;
  assign T_2379_addr_beat = 3'h0;
  assign T_2379_addr_block = xact_addr_block;
  assign T_2379_client_xact_id = xact_vol_ir_client_xact_id;
  assign T_2379_voluntary = 1'h1;
  assign T_2379_r_type = xact_vol_ir_r_type;
  assign T_2379_data = 64'h0;
  assign T_2379_client_id = xact_vol_ir_src;
  assign T_2440_addr_beat = 3'h0;
  assign T_2440_client_xact_id = T_2379_client_xact_id;
  assign T_2440_manager_xact_id = 2'h0;
  assign T_2440_is_builtin_type = 1'h1;
  assign T_2440_g_type = 4'h0;
  assign T_2440_data = 64'h0;
  assign T_2440_client_id = T_2379_client_id;
  assign GEN_0 = GEN_77;
  assign GEN_71 = 3'h1 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_72 = 3'h2 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_71;
  assign GEN_73 = 3'h3 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_72;
  assign GEN_74 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_73;
  assign GEN_75 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_74;
  assign GEN_76 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_75;
  assign GEN_77 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_76;
  assign T_2521 = GEN_0[0];
  assign GEN_1 = GEN_77;
  assign T_2522 = GEN_1[1];
  assign GEN_2 = GEN_77;
  assign T_2523 = GEN_2[2];
  assign GEN_3 = GEN_77;
  assign T_2524 = GEN_3[3];
  assign GEN_4 = GEN_77;
  assign T_2525 = GEN_4[4];
  assign GEN_5 = GEN_77;
  assign T_2526 = GEN_5[5];
  assign GEN_6 = GEN_77;
  assign T_2527 = GEN_6[6];
  assign GEN_7 = GEN_77;
  assign T_2528 = GEN_7[7];
  assign T_2532 = T_2521 ? 8'hff : 8'h0;
  assign T_2536 = T_2522 ? 8'hff : 8'h0;
  assign T_2540 = T_2523 ? 8'hff : 8'h0;
  assign T_2544 = T_2524 ? 8'hff : 8'h0;
  assign T_2548 = T_2525 ? 8'hff : 8'h0;
  assign T_2552 = T_2526 ? 8'hff : 8'h0;
  assign T_2556 = T_2527 ? 8'hff : 8'h0;
  assign T_2560 = T_2528 ? 8'hff : 8'h0;
  assign T_2561 = {T_2536,T_2532};
  assign T_2562 = {T_2544,T_2540};
  assign T_2563 = {T_2562,T_2561};
  assign T_2564 = {T_2552,T_2548};
  assign T_2565 = {T_2560,T_2556};
  assign T_2566 = {T_2565,T_2564};
  assign T_2567 = {T_2566,T_2563};
  assign T_2568 = ~ T_2567;
  assign T_2569 = T_2568 & io_inner_release_bits_data;
  assign GEN_8 = GEN_133;
  assign GEN_127 = 3'h1 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_128 = 3'h2 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_127;
  assign GEN_129 = 3'h3 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_128;
  assign GEN_130 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_129;
  assign GEN_131 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_130;
  assign GEN_132 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_131;
  assign GEN_133 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_132;
  assign T_2570 = T_2567 & GEN_8;
  assign T_2571 = T_2569 | T_2570;
  assign GEN_9 = T_2571;
  assign GEN_134 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_135 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_136 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_137 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_138 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_139 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_140 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_141 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_10 = 8'hff;
  assign GEN_142 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_0;
  assign GEN_143 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_1;
  assign GEN_144 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_2;
  assign GEN_145 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_3;
  assign GEN_146 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_4;
  assign GEN_147 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_5;
  assign GEN_148 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_6;
  assign GEN_149 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_7;
  assign GEN_160 = T_2303 ? GEN_134 : data_buffer_0;
  assign GEN_161 = T_2303 ? GEN_135 : data_buffer_1;
  assign GEN_162 = T_2303 ? GEN_136 : data_buffer_2;
  assign GEN_163 = T_2303 ? GEN_137 : data_buffer_3;
  assign GEN_164 = T_2303 ? GEN_138 : data_buffer_4;
  assign GEN_165 = T_2303 ? GEN_139 : data_buffer_5;
  assign GEN_166 = T_2303 ? GEN_140 : data_buffer_6;
  assign GEN_167 = T_2303 ? GEN_141 : data_buffer_7;
  assign GEN_169 = T_2303 ? GEN_142 : wmask_buffer_0;
  assign GEN_170 = T_2303 ? GEN_143 : wmask_buffer_1;
  assign GEN_171 = T_2303 ? GEN_144 : wmask_buffer_2;
  assign GEN_172 = T_2303 ? GEN_145 : wmask_buffer_3;
  assign GEN_173 = T_2303 ? GEN_146 : wmask_buffer_4;
  assign GEN_174 = T_2303 ? GEN_147 : wmask_buffer_5;
  assign GEN_175 = T_2303 ? GEN_148 : wmask_buffer_6;
  assign GEN_176 = T_2303 ? GEN_149 : wmask_buffer_7;
  assign T_2604_state = 2'h2;
  assign T_2631 = T_1653 | io_alloc_irel_should;
  assign T_2647 = T_2307 & T_2310;
  assign T_2648 = pending_orel_data | T_2647;
  assign T_2651 = io_outer_release_bits_r_type == 3'h0;
  assign T_2652 = io_outer_release_bits_r_type == 3'h1;
  assign T_2653 = io_outer_release_bits_r_type == 3'h2;
  assign T_2654 = T_2651 | T_2652;
  assign T_2655 = T_2654 | T_2653;
  assign T_2656 = T_2255 & T_2655;
  assign T_2660 = T_2656 ? 8'hff : 8'h0;
  assign T_2661 = ~ T_2660;
  assign T_2663 = 8'h1 << io_outer_release_bits_addr_beat;
  assign T_2664 = ~ T_2663;
  assign T_2665 = T_2661 | T_2664;
  assign T_2666 = T_2648 & T_2665;
  assign GEN_177 = T_2631 ? T_2666 : pending_orel_data;
  assign T_2677 = T_2655 == 1'h0;
  assign T_2679 = io_outer_release_bits_addr_beat == 3'h0;
  assign T_2680 = T_2677 | T_2679;
  assign GEN_179 = T_2680 ? 1'h1 : sending_orel;
  assign T_2692 = io_outer_release_bits_addr_beat == 3'h7;
  assign T_2693 = T_2677 | T_2692;
  assign GEN_180 = T_2693 ? 1'h0 : GEN_179;
  assign GEN_181 = T_2255 ? GEN_180 : sending_orel;
  assign GEN_182 = T_2255 ? 1'h0 : pending_orel_send;
  assign T_2702 = T_2255 & io_outer_release_bits_voluntary;
  assign T_2710 = T_2702 & T_2655;
  assign T_2714 = T_2712 == 3'h7;
  assign T_2716 = T_2712 + 3'h1;
  assign T_2717 = T_2716[2:0];
  assign GEN_183 = T_2710 ? T_2717 : T_2712;
  assign T_2718 = T_2710 & T_2714;
  assign T_2719 = T_2655 ? T_2712 : 3'h0;
  assign T_2720 = T_2655 ? T_2718 : T_2702;
  assign T_2723 = io_outer_grant_bits_g_type == 4'h0;
  assign T_2724 = io_outer_grant_bits_is_builtin_type & T_2723;
  assign T_2725 = T_2241 & T_2724;
  assign T_2733_0 = 3'h5;
  assign GEN_413 = {{1'd0}, T_2733_0};
  assign T_2735 = io_outer_grant_bits_g_type == GEN_413;
  assign T_2737 = io_outer_grant_bits_is_builtin_type ? T_2735 : T_2723;
  assign T_2739 = T_2725 & T_2737;
  assign T_2743 = T_2741 == 3'h7;
  assign T_2745 = T_2741 + 3'h1;
  assign T_2746 = T_2745[2:0];
  assign GEN_184 = T_2739 ? T_2746 : T_2741;
  assign T_2747 = T_2739 & T_2743;
  assign T_2748 = T_2737 ? T_2741 : 3'h0;
  assign T_2749 = T_2737 ? T_2747 : T_2725;
  assign T_2753 = T_2749 == 1'h0;
  assign T_2754 = T_2720 & T_2753;
  assign T_2756 = T_2751 + 1'h1;
  assign T_2757 = T_2756[0:0];
  assign GEN_185 = T_2754 ? T_2757 : T_2751;
  assign T_2759 = T_2720 == 1'h0;
  assign T_2760 = T_2749 & T_2759;
  assign T_2762 = T_2751 - 1'h1;
  assign T_2763 = T_2762[0:0];
  assign GEN_186 = T_2760 ? T_2763 : GEN_185;
  assign T_2765 = T_2751 > 1'h0;
  assign T_2774 = pending_orel_data >> vol_ognt_counter_up_idx;
  assign T_2775 = T_2774[0];
  assign T_2776 = T_2655 ? T_2775 : pending_orel_send;
  assign T_2777 = T_2337 & T_2776;
  assign T_2791 = T_2604_state == 2'h2;
  assign T_2792 = T_2791 ? 3'h0 : 3'h3;
  assign T_2828_addr_beat = vol_ognt_counter_up_idx;
  assign T_2828_addr_block = xact_addr_block;
  assign T_2828_client_xact_id = 2'h0;
  assign T_2828_voluntary = 1'h1;
  assign T_2828_r_type = T_2792;
  assign T_2828_data = GEN_11;
  assign GEN_11 = GEN_193;
  assign GEN_187 = 3'h1 == vol_ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_188 = 3'h2 == vol_ognt_counter_up_idx ? data_buffer_2 : GEN_187;
  assign GEN_189 = 3'h3 == vol_ognt_counter_up_idx ? data_buffer_3 : GEN_188;
  assign GEN_190 = 3'h4 == vol_ognt_counter_up_idx ? data_buffer_4 : GEN_189;
  assign GEN_191 = 3'h5 == vol_ognt_counter_up_idx ? data_buffer_5 : GEN_190;
  assign GEN_192 = 3'h6 == vol_ognt_counter_up_idx ? data_buffer_6 : GEN_191;
  assign GEN_193 = 3'h7 == vol_ognt_counter_up_idx ? data_buffer_7 : GEN_192;
  assign T_2857 = xact_iacq_is_builtin_type == 1'h0;
  assign T_2860 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_2871_0 = 3'h3;
  assign T_2873 = io_outer_acquire_bits_a_type == T_2871_0;
  assign T_2874 = io_outer_acquire_bits_is_builtin_type & T_2873;
  assign T_2875 = T_2860 & T_2874;
  assign T_2879 = T_2877 == 3'h7;
  assign T_2881 = T_2877 + 3'h1;
  assign T_2882 = T_2881[2:0];
  assign GEN_195 = T_2875 ? T_2882 : T_2877;
  assign T_2883 = T_2875 & T_2879;
  assign T_2884 = T_2874 ? T_2877 : xact_addr_beat;
  assign T_2885 = T_2874 ? T_2883 : T_2860;
  assign T_2891 = T_2724 == 1'h0;
  assign T_2892 = T_2241 & T_2891;
  assign T_2900_0 = 3'h5;
  assign GEN_414 = {{1'd0}, T_2900_0};
  assign T_2902 = io_outer_grant_bits_g_type == GEN_414;
  assign T_2904 = io_outer_grant_bits_is_builtin_type ? T_2902 : T_2723;
  assign T_2906 = T_2892 & T_2904;
  assign T_2910 = T_2908 == 3'h7;
  assign T_2912 = T_2908 + 3'h1;
  assign T_2913 = T_2912[2:0];
  assign GEN_196 = T_2906 ? T_2913 : T_2908;
  assign T_2914 = T_2906 & T_2910;
  assign T_2915 = T_2904 ? T_2908 : xact_addr_beat;
  assign T_2916 = T_2904 ? T_2914 : T_2892;
  assign T_2920 = T_2916 == 1'h0;
  assign T_2921 = T_2885 & T_2920;
  assign T_2923 = T_2918 + 1'h1;
  assign T_2924 = T_2923[0:0];
  assign GEN_197 = T_2921 ? T_2924 : T_2918;
  assign T_2926 = T_2885 == 1'h0;
  assign T_2927 = T_2916 & T_2926;
  assign T_2929 = T_2918 - 1'h1;
  assign T_2930 = T_2929[0:0];
  assign GEN_198 = T_2927 ? T_2930 : GEN_197;
  assign T_2932 = T_2918 > 1'h0;
  assign T_2933 = state == 4'h6;
  assign T_2937 = pending_put_data >> ognt_counter_up_idx;
  assign T_2938 = T_2937[0];
  assign T_2940 = T_2938 == 1'h0;
  assign T_2949_0 = 3'h2;
  assign T_2949_1 = 3'h3;
  assign T_2949_2 = 3'h4;
  assign T_2967 = xact_allocate | T_2940;
  assign T_2968 = T_2933 & T_2967;
  assign T_2971 = xact_op_code == 5'h1;
  assign T_2972 = xact_op_code == 5'h7;
  assign T_2973 = T_2971 | T_2972;
  assign T_2974 = xact_op_code[3];
  assign T_2975 = xact_op_code == 5'h4;
  assign T_2976 = T_2974 | T_2975;
  assign T_2977 = T_2973 | T_2976;
  assign T_2978 = xact_op_code == 5'h3;
  assign T_2979 = T_2977 | T_2978;
  assign T_2980 = xact_op_code == 5'h6;
  assign T_2981 = T_2979 | T_2980;
  assign T_2984 = {xact_op_code,1'h1};
  assign T_3015_addr_block = xact_addr_block;
  assign T_3015_client_xact_id = 2'h0;
  assign T_3015_addr_beat = 3'h0;
  assign T_3015_is_builtin_type = 1'h0;
  assign T_3015_a_type = {{2'd0}, T_2981};
  assign T_3015_union = {{5'd0}, T_2984};
  assign T_3015_data = 64'h0;
  assign GEN_12 = GEN_205;
  assign GEN_199 = 3'h1 == ognt_counter_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_200 = 3'h2 == ognt_counter_up_idx ? wmask_buffer_2 : GEN_199;
  assign GEN_201 = 3'h3 == ognt_counter_up_idx ? wmask_buffer_3 : GEN_200;
  assign GEN_202 = 3'h4 == ognt_counter_up_idx ? wmask_buffer_4 : GEN_201;
  assign GEN_203 = 3'h5 == ognt_counter_up_idx ? wmask_buffer_5 : GEN_202;
  assign GEN_204 = 3'h6 == ognt_counter_up_idx ? wmask_buffer_6 : GEN_203;
  assign GEN_205 = 3'h7 == ognt_counter_up_idx ? wmask_buffer_7 : GEN_204;
  assign T_3080 = {xact_op_code,1'h0};
  assign T_3081 = {xact_addr_byte,xact_op_size};
  assign T_3082 = {T_3081,T_3080};
  assign T_3084 = {xact_op_size,xact_op_code};
  assign T_3085 = {T_3084,1'h0};
  assign T_3087 = {GEN_12,1'h0};
  assign T_3099 = T_1993 ? 6'h2 : 6'h0;
  assign T_3101 = T_1995 ? 6'h0 : T_3099;
  assign T_3103 = T_1991 ? T_3082 : {{5'd0}, T_3101};
  assign T_3105 = T_2001 ? {{2'd0}, T_3087} : T_3103;
  assign T_3107 = T_1997 ? {{2'd0}, T_3087} : T_3105;
  assign T_3109 = T_2003 ? {{3'd0}, T_3085} : T_3107;
  assign T_3111 = T_1999 ? T_3082 : T_3109;
  assign T_3140_addr_block = xact_addr_block;
  assign T_3140_client_xact_id = 2'h0;
  assign T_3140_addr_beat = ognt_counter_up_idx;
  assign T_3140_is_builtin_type = 1'h1;
  assign T_3140_a_type = xact_iacq_a_type;
  assign T_3140_union = T_3111;
  assign T_3140_data = GEN_13;
  assign GEN_13 = GEN_212;
  assign GEN_206 = 3'h1 == ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_207 = 3'h2 == ognt_counter_up_idx ? data_buffer_2 : GEN_206;
  assign GEN_208 = 3'h3 == ognt_counter_up_idx ? data_buffer_3 : GEN_207;
  assign GEN_209 = 3'h4 == ognt_counter_up_idx ? data_buffer_4 : GEN_208;
  assign GEN_210 = 3'h5 == ognt_counter_up_idx ? data_buffer_5 : GEN_209;
  assign GEN_211 = 3'h6 == ognt_counter_up_idx ? data_buffer_6 : GEN_210;
  assign GEN_212 = 3'h7 == ognt_counter_up_idx ? data_buffer_7 : GEN_211;
  assign T_3168_addr_block = T_2857 ? T_3015_addr_block : T_3140_addr_block;
  assign T_3168_client_xact_id = T_2857 ? T_3015_client_xact_id : T_3140_client_xact_id;
  assign T_3168_addr_beat = T_2857 ? T_3015_addr_beat : T_3140_addr_beat;
  assign T_3168_is_builtin_type = T_2857 ? T_3015_is_builtin_type : T_3140_is_builtin_type;
  assign T_3168_a_type = T_2857 ? T_3015_a_type : T_3140_a_type;
  assign T_3168_union = T_2857 ? T_3015_union : T_3140_union;
  assign T_3168_data = T_2857 ? T_3015_data : T_3140_data;
  assign T_3197 = T_2933 & ognt_counter_up_done;
  assign GEN_213 = T_3197 ? 4'h7 : GEN_58;
  assign GEN_214 = ognt_counter_pending ? 1'h1 : vol_ognt_counter_pending;
  assign T_3207_0 = 3'h5;
  assign T_3207_1 = 3'h4;
  assign GEN_415 = {{1'd0}, T_3207_0};
  assign T_3209 = io_outer_grant_bits_g_type == GEN_415;
  assign GEN_416 = {{1'd0}, T_3207_1};
  assign T_3210 = io_outer_grant_bits_g_type == GEN_416;
  assign T_3211 = T_3209 | T_3210;
  assign T_3213 = io_outer_grant_bits_is_builtin_type ? T_3211 : T_2723;
  assign T_3214 = T_2241 & T_3213;
  assign GEN_14 = GEN_221;
  assign GEN_215 = 3'h1 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_216 = 3'h2 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_215;
  assign GEN_217 = 3'h3 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_216;
  assign GEN_218 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_217;
  assign GEN_219 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_218;
  assign GEN_220 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_219;
  assign GEN_221 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_220;
  assign T_3215 = GEN_14[0];
  assign GEN_15 = GEN_221;
  assign T_3216 = GEN_15[1];
  assign GEN_16 = GEN_221;
  assign T_3217 = GEN_16[2];
  assign GEN_17 = GEN_221;
  assign T_3218 = GEN_17[3];
  assign GEN_18 = GEN_221;
  assign T_3219 = GEN_18[4];
  assign GEN_19 = GEN_221;
  assign T_3220 = GEN_19[5];
  assign GEN_20 = GEN_221;
  assign T_3221 = GEN_20[6];
  assign GEN_21 = GEN_221;
  assign T_3222 = GEN_21[7];
  assign T_3226 = T_3215 ? 8'hff : 8'h0;
  assign T_3230 = T_3216 ? 8'hff : 8'h0;
  assign T_3234 = T_3217 ? 8'hff : 8'h0;
  assign T_3238 = T_3218 ? 8'hff : 8'h0;
  assign T_3242 = T_3219 ? 8'hff : 8'h0;
  assign T_3246 = T_3220 ? 8'hff : 8'h0;
  assign T_3250 = T_3221 ? 8'hff : 8'h0;
  assign T_3254 = T_3222 ? 8'hff : 8'h0;
  assign T_3255 = {T_3230,T_3226};
  assign T_3256 = {T_3238,T_3234};
  assign T_3257 = {T_3256,T_3255};
  assign T_3258 = {T_3246,T_3242};
  assign T_3259 = {T_3254,T_3250};
  assign T_3260 = {T_3259,T_3258};
  assign T_3261 = {T_3260,T_3257};
  assign T_3262 = ~ T_3261;
  assign T_3263 = T_3262 & io_outer_grant_bits_data;
  assign GEN_22 = GEN_277;
  assign GEN_271 = 3'h1 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_272 = 3'h2 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_271;
  assign GEN_273 = 3'h3 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_272;
  assign GEN_274 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_273;
  assign GEN_275 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_274;
  assign GEN_276 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_275;
  assign GEN_277 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_276;
  assign T_3264 = T_3261 & GEN_22;
  assign T_3265 = T_3263 | T_3264;
  assign GEN_23 = T_3265;
  assign GEN_278 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_160;
  assign GEN_279 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_161;
  assign GEN_280 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_162;
  assign GEN_281 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_163;
  assign GEN_282 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_164;
  assign GEN_283 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_165;
  assign GEN_284 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_166;
  assign GEN_285 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_167;
  assign GEN_24 = 8'hff;
  assign GEN_286 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_169;
  assign GEN_287 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_170;
  assign GEN_288 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_171;
  assign GEN_289 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_172;
  assign GEN_290 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_173;
  assign GEN_291 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_174;
  assign GEN_292 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_175;
  assign GEN_293 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_176;
  assign GEN_304 = T_3214 ? GEN_278 : GEN_160;
  assign GEN_305 = T_3214 ? GEN_279 : GEN_161;
  assign GEN_306 = T_3214 ? GEN_280 : GEN_162;
  assign GEN_307 = T_3214 ? GEN_281 : GEN_163;
  assign GEN_308 = T_3214 ? GEN_282 : GEN_164;
  assign GEN_309 = T_3214 ? GEN_283 : GEN_165;
  assign GEN_310 = T_3214 ? GEN_284 : GEN_166;
  assign GEN_311 = T_3214 ? GEN_285 : GEN_167;
  assign GEN_313 = T_3214 ? GEN_286 : GEN_169;
  assign GEN_314 = T_3214 ? GEN_287 : GEN_170;
  assign GEN_315 = T_3214 ? GEN_288 : GEN_171;
  assign GEN_316 = T_3214 ? GEN_289 : GEN_172;
  assign GEN_317 = T_3214 ? GEN_290 : GEN_173;
  assign GEN_318 = T_3214 ? GEN_291 : GEN_174;
  assign GEN_319 = T_3214 ? GEN_292 : GEN_175;
  assign GEN_320 = T_3214 ? GEN_293 : GEN_176;
  assign T_3268 = scoreboard_3 | ognt_counter_pending;
  assign T_3269 = T_3268 | vol_ognt_counter_pending;
  assign T_3281 = T_2179 == 1'h0;
  assign T_3283 = T_2175 & T_3281;
  assign T_3291_0 = 3'h5;
  assign GEN_417 = {{1'd0}, T_3291_0};
  assign T_3293 = io_inner_grant_bits_g_type == GEN_417;
  assign T_3295 = io_inner_grant_bits_is_builtin_type ? T_3293 : T_2178;
  assign T_3297 = T_3283 & T_3295;
  assign T_3301 = T_3299 == 3'h7;
  assign T_3303 = T_3299 + 3'h1;
  assign T_3304 = T_3303[2:0];
  assign GEN_321 = T_3297 ? T_3304 : T_3299;
  assign T_3305 = T_3297 & T_3301;
  assign T_3306 = T_3295 ? T_3299 : 3'h0;
  assign T_3307 = T_3295 ? T_3305 : T_3283;
  assign T_3308 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3326 = T_3308 == 1'h0;
  assign T_3327 = T_3307 & T_3326;
  assign T_3329 = T_3324 + 1'h1;
  assign T_3330 = T_3329[0:0];
  assign GEN_323 = T_3327 ? T_3330 : T_3324;
  assign T_3332 = T_3307 == 1'h0;
  assign T_3333 = T_3308 & T_3332;
  assign T_3335 = T_3324 - 1'h1;
  assign T_3336 = T_3335[0:0];
  assign GEN_324 = T_3333 ? T_3336 : GEN_323;
  assign T_3338 = T_3324 > 1'h0;
  assign T_3343 = T_1798 == 1'h0;
  assign T_3360 = pending_ignt_data | T_2647;
  assign T_3370_0 = 3'h5;
  assign T_3370_1 = 3'h4;
  assign GEN_418 = {{1'd0}, T_3370_0};
  assign T_3372 = io_outer_grant_bits_g_type == GEN_418;
  assign GEN_419 = {{1'd0}, T_3370_1};
  assign T_3373 = io_outer_grant_bits_g_type == GEN_419;
  assign T_3374 = T_3372 | T_3373;
  assign T_3376 = io_outer_grant_bits_is_builtin_type ? T_3374 : T_2723;
  assign T_3377 = T_2241 & T_3376;
  assign T_3382 = T_3377 ? 8'hff : 8'h0;
  assign T_3384 = 8'h1 << io_outer_grant_bits_addr_beat;
  assign T_3385 = T_3382 & T_3384;
  assign T_3386 = T_3360 | T_3385;
  assign GEN_327 = T_3343 ? T_3386 : GEN_45;
  assign T_3389 = state == 4'h1;
  assign T_3390 = T_1611 | T_3389;
  assign T_3393 = T_3390 | scoreboard_0;
  assign T_3395 = T_3393 == 1'h0;
  assign T_3412 = 3'h6 == ignt_q_io_deq_bits_a_type;
  assign T_3413 = T_3412 ? 3'h1 : 3'h3;
  assign T_3414 = 3'h5 == ignt_q_io_deq_bits_a_type;
  assign T_3415 = T_3414 ? 3'h1 : T_3413;
  assign T_3416 = 3'h4 == ignt_q_io_deq_bits_a_type;
  assign T_3417 = T_3416 ? 3'h4 : T_3415;
  assign T_3418 = 3'h3 == ignt_q_io_deq_bits_a_type;
  assign T_3419 = T_3418 ? 3'h3 : T_3417;
  assign T_3420 = 3'h2 == ignt_q_io_deq_bits_a_type;
  assign T_3421 = T_3420 ? 3'h3 : T_3419;
  assign T_3422 = 3'h1 == ignt_q_io_deq_bits_a_type;
  assign T_3423 = T_3422 ? 3'h5 : T_3421;
  assign T_3424 = 3'h0 == ignt_q_io_deq_bits_a_type;
  assign T_3425 = T_3424 ? 3'h4 : T_3423;
  assign T_3426 = ignt_q_io_deq_bits_is_builtin_type ? T_3425 : 3'h0;
  assign T_3455_addr_beat = ignt_q_io_deq_bits_addr_beat;
  assign T_3455_client_xact_id = ignt_q_io_deq_bits_client_xact_id;
  assign T_3455_manager_xact_id = 2'h1;
  assign T_3455_is_builtin_type = ignt_q_io_deq_bits_is_builtin_type;
  assign T_3455_g_type = {{1'd0}, T_3426};
  assign T_3455_data = GEN_25;
  assign T_3455_client_id = ignt_q_io_deq_bits_client_id;
  assign GEN_25 = GEN_334;
  assign GEN_328 = 3'h1 == ignt_data_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_329 = 3'h2 == ignt_data_idx ? data_buffer_2 : GEN_328;
  assign GEN_330 = 3'h3 == ignt_data_idx ? data_buffer_3 : GEN_329;
  assign GEN_331 = 3'h4 == ignt_data_idx ? data_buffer_4 : GEN_330;
  assign GEN_332 = 3'h5 == ignt_data_idx ? data_buffer_5 : GEN_331;
  assign GEN_333 = 3'h6 == ignt_data_idx ? data_buffer_6 : GEN_332;
  assign GEN_334 = 3'h7 == ignt_data_idx ? data_buffer_7 : GEN_333;
  assign T_3491_0 = 3'h5;
  assign GEN_420 = {{1'd0}, T_3491_0};
  assign T_3493 = io_inner_grant_bits_g_type == GEN_420;
  assign T_3495 = io_inner_grant_bits_is_builtin_type ? T_3493 : T_2178;
  assign T_3497 = T_2175 & T_3495;
  assign T_3501 = T_3499 == 3'h7;
  assign T_3503 = T_3499 + 3'h1;
  assign T_3504 = T_3503[2:0];
  assign GEN_335 = T_3497 ? T_3504 : T_3499;
  assign T_3505 = T_3497 & T_3501;
  assign T_3506 = T_3495 ? T_3499 : ignt_q_io_deq_bits_addr_beat;
  assign T_3507 = T_3495 ? T_3505 : T_2175;
  assign T_3512 = T_2337 & scoreboard_6;
  assign T_3514 = T_3269 == 1'h0;
  assign T_3522_0 = 3'h5;
  assign T_3522_1 = 3'h4;
  assign GEN_421 = {{1'd0}, T_3522_0};
  assign T_3524 = io_inner_grant_bits_g_type == GEN_421;
  assign GEN_422 = {{1'd0}, T_3522_1};
  assign T_3525 = io_inner_grant_bits_g_type == GEN_422;
  assign T_3526 = T_3524 | T_3525;
  assign T_3528 = io_inner_grant_bits_is_builtin_type ? T_3526 : T_2178;
  assign T_3529 = pending_ignt_data >> ignt_data_idx;
  assign T_3530 = T_3529[0];
  assign T_3532 = T_3528 ? T_3530 : T_3395;
  assign T_3533 = T_3514 & T_3532;
  assign GEN_338 = T_3512 ? T_3533 : T_2347;
  assign GEN_339 = T_2250 ? ignt_data_done : 1'h0;
  assign GEN_340 = T_2250 ? ignt_data_idx : T_2440_addr_beat;
  assign GEN_341 = T_2250 ? T_3455_client_xact_id : T_2440_client_xact_id;
  assign GEN_342 = T_2250 ? T_3455_manager_xact_id : T_2440_manager_xact_id;
  assign GEN_343 = T_2250 ? T_3455_is_builtin_type : T_2440_is_builtin_type;
  assign GEN_344 = T_2250 ? T_3455_g_type : T_2440_g_type;
  assign GEN_345 = T_2250 ? T_3455_data : T_2440_data;
  assign GEN_346 = T_2250 ? T_3455_client_id : T_2440_client_id;
  assign GEN_349 = T_2250 ? GEN_338 : T_2347;
  assign T_3540 = ~ io_incoherent_0;
  assign GEN_350 = T_1798 ? {{1'd0}, T_3540} : T_2079;
  assign T_3551 = T_1767 & io_inner_acquire_valid;
  assign T_3552 = T_1798 | T_3551;
  assign T_3562_0 = 3'h2;
  assign T_3562_1 = 3'h3;
  assign T_3562_2 = 3'h4;
  assign T_3564 = io_inner_acquire_bits_a_type == T_3562_0;
  assign T_3565 = io_inner_acquire_bits_a_type == T_3562_1;
  assign T_3566 = io_inner_acquire_bits_a_type == T_3562_2;
  assign T_3567 = T_3564 | T_3565;
  assign T_3568 = T_3567 | T_3566;
  assign T_3569 = io_inner_acquire_bits_is_builtin_type & T_3568;
  assign T_3570 = T_1612 & T_3569;
  assign T_3571 = T_3570 & T_3552;
  assign T_3573 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3574 = io_inner_acquire_bits_is_builtin_type & T_3573;
  assign T_3603 = T_1921 | T_1918;
  assign T_3604 = io_inner_acquire_bits_union[8:1];
  assign T_3606 = T_3603 ? T_3604 : 8'h0;
  assign T_3607 = T_3574 ? 8'hff : T_3606;
  assign T_3608 = T_3607[0];
  assign T_3609 = T_3607[1];
  assign T_3610 = T_3607[2];
  assign T_3611 = T_3607[3];
  assign T_3612 = T_3607[4];
  assign T_3613 = T_3607[5];
  assign T_3614 = T_3607[6];
  assign T_3615 = T_3607[7];
  assign T_3619 = T_3608 ? 8'hff : 8'h0;
  assign T_3623 = T_3609 ? 8'hff : 8'h0;
  assign T_3627 = T_3610 ? 8'hff : 8'h0;
  assign T_3631 = T_3611 ? 8'hff : 8'h0;
  assign T_3635 = T_3612 ? 8'hff : 8'h0;
  assign T_3639 = T_3613 ? 8'hff : 8'h0;
  assign T_3643 = T_3614 ? 8'hff : 8'h0;
  assign T_3647 = T_3615 ? 8'hff : 8'h0;
  assign T_3648 = {T_3623,T_3619};
  assign T_3649 = {T_3631,T_3627};
  assign T_3650 = {T_3649,T_3648};
  assign T_3651 = {T_3639,T_3635};
  assign T_3652 = {T_3647,T_3643};
  assign T_3653 = {T_3652,T_3651};
  assign T_3654 = {T_3653,T_3650};
  assign T_3655 = ~ T_3654;
  assign GEN_26 = GEN_357;
  assign GEN_351 = 3'h1 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_352 = 3'h2 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_351;
  assign GEN_353 = 3'h3 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_352;
  assign GEN_354 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_353;
  assign GEN_355 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_354;
  assign GEN_356 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_355;
  assign GEN_357 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_356;
  assign T_3656 = T_3655 & GEN_26;
  assign T_3657 = T_3654 & io_inner_acquire_bits_data;
  assign T_3658 = T_3656 | T_3657;
  assign GEN_27 = T_3658;
  assign GEN_358 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_304;
  assign GEN_359 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_305;
  assign GEN_360 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_306;
  assign GEN_361 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_307;
  assign GEN_362 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_308;
  assign GEN_363 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_309;
  assign GEN_364 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_310;
  assign GEN_365 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_311;
  assign GEN_28 = GEN_372;
  assign GEN_366 = 3'h1 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_367 = 3'h2 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_366;
  assign GEN_368 = 3'h3 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_367;
  assign GEN_369 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_368;
  assign GEN_370 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_369;
  assign GEN_371 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_370;
  assign GEN_372 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_371;
  assign T_3695 = T_3607 | GEN_28;
  assign GEN_29 = T_3695;
  assign GEN_373 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_313;
  assign GEN_374 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_314;
  assign GEN_375 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_315;
  assign GEN_376 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_316;
  assign GEN_377 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_317;
  assign GEN_378 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_318;
  assign GEN_379 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_319;
  assign GEN_380 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_320;
  assign GEN_383 = T_3571 ? GEN_358 : GEN_304;
  assign GEN_384 = T_3571 ? GEN_359 : GEN_305;
  assign GEN_385 = T_3571 ? GEN_360 : GEN_306;
  assign GEN_386 = T_3571 ? GEN_361 : GEN_307;
  assign GEN_387 = T_3571 ? GEN_362 : GEN_308;
  assign GEN_388 = T_3571 ? GEN_363 : GEN_309;
  assign GEN_389 = T_3571 ? GEN_364 : GEN_310;
  assign GEN_390 = T_3571 ? GEN_365 : GEN_311;
  assign GEN_393 = T_3571 ? GEN_373 : GEN_313;
  assign GEN_394 = T_3571 ? GEN_374 : GEN_314;
  assign GEN_395 = T_3571 ? GEN_375 : GEN_315;
  assign GEN_396 = T_3571 ? GEN_376 : GEN_316;
  assign GEN_397 = T_3571 ? GEN_377 : GEN_317;
  assign GEN_398 = T_3571 ? GEN_378 : GEN_318;
  assign GEN_399 = T_3571 ? GEN_379 : GEN_319;
  assign GEN_400 = T_3571 ? GEN_380 : GEN_320;
  assign T_3698 = scoreboard_0 | T_2343;
  assign T_3699 = T_3698 | vol_ignt_counter_pending;
  assign T_3700 = T_3699 | scoreboard_3;
  assign T_3701 = T_3700 | vol_ognt_counter_pending;
  assign T_3702 = T_3701 | ognt_counter_pending;
  assign T_3703 = T_3702 | scoreboard_6;
  assign T_3704 = T_3703 | ifin_counter_pending;
  assign T_3706 = T_3704 == 1'h0;
  assign T_3708 = T_2337 & all_pending_done;
  assign GEN_401 = T_3708 ? 4'h0 : GEN_213;
  assign GEN_402 = T_3708 ? 8'h0 : GEN_393;
  assign GEN_403 = T_3708 ? 8'h0 : GEN_394;
  assign GEN_404 = T_3708 ? 8'h0 : GEN_395;
  assign GEN_405 = T_3708 ? 8'h0 : GEN_396;
  assign GEN_406 = T_3708 ? 8'h0 : GEN_397;
  assign GEN_407 = T_3708 ? 8'h0 : GEN_398;
  assign GEN_408 = T_3708 ? 8'h0 : GEN_399;
  assign GEN_409 = T_3708 ? 8'h0 : GEN_400;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_121[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_122[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  state = GEN_32[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  xact_addr_block = GEN_33[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  xact_allocate = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  xact_amo_shift_bytes = GEN_42[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  xact_op_code = GEN_43[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  xact_addr_byte = GEN_47[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_78 = {1{$random}};
  xact_op_size = GEN_78[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_79 = {1{$random}};
  xact_vol_ir_r_type = GEN_79[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_80 = {1{$random}};
  xact_vol_ir_src = GEN_80[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_81 = {1{$random}};
  xact_vol_ir_client_xact_id = GEN_81[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_82 = {1{$random}};
  pending_irel_data = GEN_82[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_83 = {1{$random}};
  pending_put_data = GEN_83[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_84 = {1{$random}};
  pending_ignt_data = GEN_84[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {1{$random}};
  pending_iprbs = GEN_85[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  pending_orel_send = GEN_86[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_87 = {1{$random}};
  pending_orel_data = GEN_87[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  sending_orel = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {2{$random}};
  data_buffer_0 = GEN_89[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {2{$random}};
  data_buffer_1 = GEN_90[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {2{$random}};
  data_buffer_2 = GEN_91[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_92 = {2{$random}};
  data_buffer_3 = GEN_92[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_93 = {2{$random}};
  data_buffer_4 = GEN_93[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_94 = {2{$random}};
  data_buffer_5 = GEN_94[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_95 = {2{$random}};
  data_buffer_6 = GEN_95[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_96 = {2{$random}};
  data_buffer_7 = GEN_96[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_97 = {1{$random}};
  wmask_buffer_0 = GEN_97[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_98 = {1{$random}};
  wmask_buffer_1 = GEN_98[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_99 = {1{$random}};
  wmask_buffer_2 = GEN_99[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {1{$random}};
  wmask_buffer_3 = GEN_100[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_101 = {1{$random}};
  wmask_buffer_4 = GEN_101[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_102 = {1{$random}};
  wmask_buffer_5 = GEN_102[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_103 = {1{$random}};
  wmask_buffer_6 = GEN_103[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_104 = {1{$random}};
  wmask_buffer_7 = GEN_104[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_105 = {1{$random}};
  T_2091 = GEN_105[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_106 = {1{$random}};
  T_2115 = GEN_106[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_107 = {1{$random}};
  T_2125 = GEN_107[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_108 = {1{$random}};
  T_2166 = GEN_108[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_109 = {1{$random}};
  T_2197 = GEN_109[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_110 = {1{$random}};
  T_2207 = GEN_110[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_111 = {1{$random}};
  T_2712 = GEN_111[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {1{$random}};
  T_2741 = GEN_112[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_113 = {1{$random}};
  T_2751 = GEN_113[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_114 = {1{$random}};
  T_2877 = GEN_114[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  T_2908 = GEN_115[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_116 = {1{$random}};
  T_2918 = GEN_116[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_117 = {1{$random}};
  T_3299 = GEN_117[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_118 = {1{$random}};
  T_3314 = GEN_118[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  T_3324 = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  T_3499 = GEN_120[2:0];
  `endif
  GEN_121 = {1{$random}};
  GEN_122 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_3708) begin
        state <= 4'h0;
      end else begin
        if(T_3197) begin
          state <= 4'h7;
        end else begin
          if(T_2224) begin
            state <= 4'h7;
          end else begin
            if(T_2146) begin
              if(T_2055) begin
                state <= 4'h6;
              end else begin
                state <= 4'h7;
              end
            end else begin
              if(T_1798) begin
                state <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      xact_addr_block <= 26'h0;
    end else begin
      if(T_2224) begin
        xact_addr_block <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1798) begin
          xact_addr_block <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_allocate <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_amo_shift_bytes <= T_1915;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        if(T_1922) begin
          xact_op_code <= 5'h1;
        end else begin
          xact_op_code <= T_1923;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_addr_byte <= T_1925;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_op_size <= T_1926;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_r_type <= io_inner_release_bits_r_type;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_src <= io_inner_release_bits_client_id;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_client_xact_id <= io_inner_release_bits_client_xact_id;
          end
        end
      end
    end
    if(reset) begin
      pending_irel_data <= 8'h0;
    end else begin
      if(T_2277) begin
        if(T_2316) begin
          pending_irel_data <= T_2333;
        end else begin
          if(T_2289) begin
            if(T_2111) begin
              pending_irel_data <= T_2312;
            end else begin
              pending_irel_data <= 8'h0;
            end
          end else begin
            if(T_2224) begin
              pending_irel_data <= 8'hff;
            end
          end
        end
      end else begin
        if(T_2224) begin
          pending_irel_data <= 8'hff;
        end
      end
    end
    if(reset) begin
      pending_put_data <= 8'h0;
    end else begin
      if(T_1798) begin
        if(T_1921) begin
          pending_put_data <= T_1956;
        end else begin
          pending_put_data <= 8'h0;
        end
      end else begin
        if(T_1852) begin
          pending_put_data <= T_1907;
        end
      end
    end
    if(reset) begin
      pending_ignt_data <= 8'h0;
    end else begin
      if(T_3343) begin
        pending_ignt_data <= T_3386;
      end else begin
        if(T_1798) begin
          pending_ignt_data <= 8'h0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      pending_iprbs <= GEN_350[0];
    end
    if(reset) begin
      pending_orel_send <= 1'h0;
    end else begin
      if(T_2255) begin
        pending_orel_send <= 1'h0;
      end
    end
    if(reset) begin
      pending_orel_data <= 8'h0;
    end else begin
      if(T_2631) begin
        pending_orel_data <= T_2666;
      end
    end
    if(reset) begin
      sending_orel <= 1'h0;
    end else begin
      if(T_2255) begin
        if(T_2693) begin
          sending_orel <= 1'h0;
        end else begin
          if(T_2680) begin
            sending_orel <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1691_0;
    end else begin
      if(T_3571) begin
        if(3'h0 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h0 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h0 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1691_1;
    end else begin
      if(T_3571) begin
        if(3'h1 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h1 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h1 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1691_2;
    end else begin
      if(T_3571) begin
        if(3'h2 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h2 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h2 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1691_3;
    end else begin
      if(T_3571) begin
        if(3'h3 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h3 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h3 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1691_4;
    end else begin
      if(T_3571) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1691_5;
    end else begin
      if(T_3571) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1691_6;
    end else begin
      if(T_3571) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1691_7;
    end else begin
      if(T_3571) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1709_0;
    end else begin
      if(T_3708) begin
        wmask_buffer_0 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h0 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h0 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h0 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_0 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_0 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1709_1;
    end else begin
      if(T_3708) begin
        wmask_buffer_1 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h1 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h1 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h1 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_1 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_1 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1709_2;
    end else begin
      if(T_3708) begin
        wmask_buffer_2 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h2 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h2 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h2 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_2 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_2 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1709_3;
    end else begin
      if(T_3708) begin
        wmask_buffer_3 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h3 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h3 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h3 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_3 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_3 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1709_4;
    end else begin
      if(T_3708) begin
        wmask_buffer_4 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h4 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h4 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_4 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_4 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1709_5;
    end else begin
      if(T_3708) begin
        wmask_buffer_5 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h5 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h5 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_5 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_5 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1709_6;
    end else begin
      if(T_3708) begin
        wmask_buffer_6 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h6 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h6 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_6 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_6 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1709_7;
    end else begin
      if(T_3708) begin
        wmask_buffer_7 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h7 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h7 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_7 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_7 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_2091 <= 3'h0;
    end
    if(reset) begin
      T_2115 <= 3'h0;
    end else begin
      if(T_2113) begin
        T_2115 <= T_2120;
      end
    end
    if(reset) begin
      T_2125 <= 1'h0;
    end else begin
      if(T_2134) begin
        T_2125 <= T_2137;
      end else begin
        if(T_2128) begin
          T_2125 <= T_2131;
        end
      end
    end
    if(reset) begin
      T_2166 <= 3'h0;
    end else begin
      if(T_2164) begin
        T_2166 <= T_2171;
      end
    end
    if(reset) begin
      T_2197 <= 3'h0;
    end else begin
      if(T_2195) begin
        T_2197 <= T_2202;
      end
    end
    if(reset) begin
      T_2207 <= 1'h0;
    end else begin
      if(T_2216) begin
        T_2207 <= T_2219;
      end else begin
        if(T_2210) begin
          T_2207 <= T_2213;
        end
      end
    end
    if(reset) begin
      T_2712 <= 3'h0;
    end else begin
      if(T_2710) begin
        T_2712 <= T_2717;
      end
    end
    if(reset) begin
      T_2741 <= 3'h0;
    end else begin
      if(T_2739) begin
        T_2741 <= T_2746;
      end
    end
    if(reset) begin
      T_2751 <= 1'h0;
    end else begin
      if(T_2760) begin
        T_2751 <= T_2763;
      end else begin
        if(T_2754) begin
          T_2751 <= T_2757;
        end
      end
    end
    if(reset) begin
      T_2877 <= 3'h0;
    end else begin
      if(T_2875) begin
        T_2877 <= T_2882;
      end
    end
    if(reset) begin
      T_2908 <= 3'h0;
    end else begin
      if(T_2906) begin
        T_2908 <= T_2913;
      end
    end
    if(reset) begin
      T_2918 <= 1'h0;
    end else begin
      if(T_2927) begin
        T_2918 <= T_2930;
      end else begin
        if(T_2921) begin
          T_2918 <= T_2924;
        end
      end
    end
    if(reset) begin
      T_3299 <= 3'h0;
    end else begin
      if(T_3297) begin
        T_3299 <= T_3304;
      end
    end
    if(reset) begin
      T_3314 <= 3'h0;
    end
    if(reset) begin
      T_3324 <= 1'h0;
    end else begin
      if(T_3333) begin
        T_3324 <= T_3336;
      end else begin
        if(T_3327) begin
          T_3324 <= T_3330;
        end
      end
    end
    if(reset) begin
      T_3499 <= 3'h0;
    end else begin
      if(T_3497) begin
        T_3499 <= T_3504;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1652) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:98 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1652) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1666) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1677) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:105 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1677) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BufferedBroadcastAcquireTracker_1(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input   io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output  io_inner_grant_bits_client_xact_id,
  output [1:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [1:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input   io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [1:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should,
  output  io_alloc_idle,
  output [25:0] io_alloc_addr_block
);
  wire  all_pending_done;
  reg [3:0] state;
  reg [31:0] GEN_32;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_33;
  reg  xact_allocate;
  reg [31:0] GEN_41;
  reg [4:0] xact_amo_shift_bytes;
  reg [31:0] GEN_42;
  reg [4:0] xact_op_code;
  reg [31:0] GEN_43;
  reg [2:0] xact_addr_byte;
  reg [31:0] GEN_47;
  reg [1:0] xact_op_size;
  reg [31:0] GEN_78;
  wire [2:0] xact_addr_beat;
  wire  xact_iacq_client_xact_id;
  wire [2:0] xact_iacq_addr_beat;
  wire  xact_iacq_client_id;
  wire  xact_iacq_is_builtin_type;
  wire [2:0] xact_iacq_a_type;
  reg [2:0] xact_vol_ir_r_type;
  reg [31:0] GEN_79;
  reg  xact_vol_ir_src;
  reg [31:0] GEN_80;
  reg  xact_vol_ir_client_xact_id;
  reg [31:0] GEN_81;
  reg [7:0] pending_irel_data;
  reg [31:0] GEN_82;
  wire  vol_ignt_counter_pending;
  wire [2:0] vol_ignt_counter_up_idx;
  wire  vol_ignt_counter_up_done;
  wire [2:0] vol_ignt_counter_down_idx;
  wire  vol_ignt_counter_down_done;
  wire  scoreboard_6;
  wire [2:0] ignt_data_idx;
  wire  ignt_data_done;
  wire  ifin_counter_pending;
  wire [2:0] ifin_counter_up_idx;
  wire  ifin_counter_up_done;
  wire [2:0] ifin_counter_down_idx;
  wire  ifin_counter_down_done;
  reg [7:0] pending_put_data;
  reg [31:0] GEN_83;
  reg [7:0] pending_ignt_data;
  reg [31:0] GEN_84;
  wire  ognt_counter_pending;
  wire [2:0] ognt_counter_up_idx;
  wire  ognt_counter_up_done;
  wire [2:0] ognt_counter_down_idx;
  wire  ognt_counter_down_done;
  reg  pending_iprbs;
  reg [31:0] GEN_85;
  reg  pending_orel_send;
  reg [31:0] GEN_86;
  reg [7:0] pending_orel_data;
  reg [31:0] GEN_87;
  wire  vol_ognt_counter_pending;
  wire [2:0] vol_ognt_counter_up_idx;
  wire  vol_ognt_counter_up_done;
  wire [2:0] vol_ognt_counter_down_idx;
  wire  vol_ognt_counter_down_done;
  wire  T_170;
  wire  T_171;
  wire  scoreboard_3;
  reg  sending_orel;
  reg [31:0] GEN_88;
  wire  T_195_sharers;
  wire [1:0] T_241_state;
  wire  coh_inner_sharers;
  wire [1:0] coh_outer_state;
  wire  T_1611;
  wire  T_1612;
  wire  T_1613;
  wire  T_1614;
  wire [2:0] T_1623_0;
  wire  T_1625;
  wire  T_1626;
  wire  T_1627;
  wire [2:0] T_1636_0;
  wire  T_1638;
  wire  T_1639;
  wire  T_1641;
  wire  T_1643;
  wire  T_1644;
  wire  T_1646;
  wire  T_1647;
  wire  T_1649;
  wire  T_1650;
  wire  T_1652;
  wire  T_1653;
  wire  T_1654;
  wire  T_1656;
  wire  T_1658;
  wire  T_1659;
  wire  T_1660;
  wire  T_1661;
  wire  T_1663;
  wire  T_1664;
  wire  T_1666;
  wire  T_1670;
  wire  T_1671;
  wire  T_1672;
  wire  T_1674;
  wire  T_1675;
  wire  T_1677;
  wire [63:0] T_1691_0;
  wire [63:0] T_1691_1;
  wire [63:0] T_1691_2;
  wire [63:0] T_1691_3;
  wire [63:0] T_1691_4;
  wire [63:0] T_1691_5;
  wire [63:0] T_1691_6;
  wire [63:0] T_1691_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_89;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_90;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_91;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_92;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_93;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_94;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_95;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_96;
  wire [7:0] T_1709_0;
  wire [7:0] T_1709_1;
  wire [7:0] T_1709_2;
  wire [7:0] T_1709_3;
  wire [7:0] T_1709_4;
  wire [7:0] T_1709_5;
  wire [7:0] T_1709_6;
  wire [7:0] T_1709_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_97;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_98;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_99;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_100;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_101;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_102;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_103;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_104;
  wire [7:0] T_1714;
  wire  T_1716;
  wire [7:0] T_1717;
  wire  T_1719;
  wire [7:0] T_1720;
  wire  T_1722;
  wire [7:0] T_1723;
  wire  T_1725;
  wire [7:0] T_1726;
  wire  T_1728;
  wire [7:0] T_1729;
  wire  T_1731;
  wire [7:0] T_1732;
  wire  T_1734;
  wire [7:0] T_1735;
  wire  T_1737;
  wire  data_valid_0;
  wire  data_valid_1;
  wire  data_valid_2;
  wire  data_valid_3;
  wire  data_valid_4;
  wire  data_valid_5;
  wire  data_valid_6;
  wire  data_valid_7;
  wire  T_1748;
  wire  T_1749;
  wire  T_1751;
  wire  T_1752;
  wire  T_1754;
  wire  T_1755;
  wire  T_1764;
  wire  T_1765;
  wire  T_1766;
  wire  T_1767;
  wire  T_1768;
  wire  T_1769;
  wire  ignt_q_clk;
  wire  ignt_q_reset;
  wire  ignt_q_io_enq_ready;
  wire  ignt_q_io_enq_valid;
  wire  ignt_q_io_enq_bits_client_xact_id;
  wire [2:0] ignt_q_io_enq_bits_addr_beat;
  wire  ignt_q_io_enq_bits_client_id;
  wire  ignt_q_io_enq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_enq_bits_a_type;
  wire  ignt_q_io_deq_ready;
  wire  ignt_q_io_deq_valid;
  wire  ignt_q_io_deq_bits_client_xact_id;
  wire [2:0] ignt_q_io_deq_bits_addr_beat;
  wire  ignt_q_io_deq_bits_client_id;
  wire  ignt_q_io_deq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_deq_bits_a_type;
  wire [1:0] ignt_q_io_count;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [2:0] T_1812_0;
  wire  T_1814;
  wire  T_1815;
  wire  T_1817;
  wire  T_1820;
  wire  T_1821;
  wire  T_1822;
  wire  T_1823_client_xact_id;
  wire [2:0] T_1823_addr_beat;
  wire  T_1823_client_id;
  wire  T_1823_is_builtin_type;
  wire [2:0] T_1823_a_type;
  wire  T_1850;
  wire  T_1852;
  wire [2:0] T_1862_0;
  wire [2:0] T_1862_1;
  wire [2:0] T_1862_2;
  wire  T_1864;
  wire  T_1865;
  wire  T_1866;
  wire  T_1867;
  wire  T_1868;
  wire  T_1869;
  wire  T_1870;
  wire [7:0] T_1874;
  wire [7:0] T_1875;
  wire [7:0] T_1877;
  wire [7:0] T_1878;
  wire [7:0] T_1879;
  wire [7:0] T_1880;
  wire [2:0] T_1890_0;
  wire  T_1892;
  wire  T_1893;
  wire  T_1894;
  wire  T_1897;
  wire [7:0] T_1906;
  wire [7:0] T_1907;
  wire [7:0] GEN_34;
  wire [4:0] T_1915;
  wire  T_1917;
  wire  T_1918;
  wire  T_1920;
  wire  T_1921;
  wire  T_1922;
  wire [4:0] T_1923;
  wire [4:0] T_1924;
  wire [2:0] T_1925;
  wire [1:0] T_1926;
  wire [2:0] T_1939_0;
  wire [2:0] T_1939_1;
  wire [2:0] T_1939_2;
  wire  T_1941;
  wire  T_1942;
  wire  T_1943;
  wire  T_1944;
  wire  T_1945;
  wire  T_1946;
  wire  T_1947;
  wire [7:0] T_1951;
  wire [7:0] T_1952;
  wire [7:0] T_1956;
  wire [7:0] T_1958;
  wire [25:0] GEN_35;
  wire  GEN_36;
  wire [4:0] GEN_37;
  wire [4:0] GEN_38;
  wire [2:0] GEN_39;
  wire [1:0] GEN_40;
  wire [7:0] GEN_44;
  wire [7:0] GEN_45;
  wire [3:0] GEN_46;
  wire  scoreboard_0;
  wire [2:0] T_1976_0;
  wire  T_1978;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire [7:0] T_1982;
  wire  skip_outer_acquire;
  wire  T_1991;
  wire [1:0] T_1992;
  wire  T_1993;
  wire [1:0] T_1994;
  wire  T_1995;
  wire [1:0] T_1996;
  wire  T_1997;
  wire [1:0] T_1998;
  wire  T_1999;
  wire [1:0] T_2000;
  wire  T_2001;
  wire [1:0] T_2002;
  wire  T_2003;
  wire [1:0] T_2004;
  wire [1:0] T_2005;
  wire [25:0] T_2030_addr_block;
  wire [1:0] T_2030_p_type;
  wire  T_2030_client_id;
  wire  T_2055;
  wire [3:0] T_2056;
  wire  T_2065_pending;
  wire [2:0] T_2065_up_idx;
  wire  T_2065_up_done;
  wire [2:0] T_2065_down_idx;
  wire  T_2065_down_done;
  wire  T_2073;
  wire  T_2074;
  wire [1:0] T_2076;
  wire [1:0] T_2077;
  wire [1:0] GEN_410;
  wire [1:0] T_2078;
  wire [1:0] GEN_411;
  wire [1:0] T_2079;
  wire  T_2080;
  wire  T_2083;
  reg [2:0] T_2091;
  reg [31:0] GEN_105;
  wire  T_2100;
  wire  T_2103;
  wire  T_2104;
  wire  T_2105;
  wire  T_2107;
  wire  T_2108;
  wire  T_2109;
  wire  T_2110;
  wire  T_2111;
  wire  T_2113;
  reg [2:0] T_2115;
  reg [31:0] GEN_106;
  wire  T_2117;
  wire [3:0] T_2119;
  wire [2:0] T_2120;
  wire [2:0] GEN_48;
  wire  T_2121;
  wire [2:0] T_2122;
  wire  T_2123;
  reg  T_2125;
  reg [31:0] GEN_107;
  wire  T_2127;
  wire  T_2128;
  wire [1:0] T_2130;
  wire  T_2131;
  wire  GEN_49;
  wire  T_2133;
  wire  T_2134;
  wire [1:0] T_2136;
  wire  T_2137;
  wire  GEN_50;
  wire  T_2139;
  wire  T_2143;
  wire  T_2145;
  wire  T_2146;
  wire [3:0] GEN_51;
  wire  T_2150;
  wire  T_2151;
  wire  T_2156;
  wire  T_2164;
  reg [2:0] T_2166;
  reg [31:0] GEN_108;
  wire  T_2168;
  wire [3:0] T_2170;
  wire [2:0] T_2171;
  wire [2:0] GEN_52;
  wire  T_2172;
  wire [2:0] T_2173;
  wire  T_2174;
  wire  T_2175;
  wire  T_2178;
  wire  T_2179;
  wire  T_2180;
  wire  T_2181;
  wire [2:0] T_2189_0;
  wire [3:0] GEN_412;
  wire  T_2191;
  wire  T_2193;
  wire  T_2195;
  reg [2:0] T_2197;
  reg [31:0] GEN_109;
  wire  T_2199;
  wire [3:0] T_2201;
  wire [2:0] T_2202;
  wire [2:0] GEN_53;
  wire  T_2203;
  wire [2:0] T_2204;
  wire  T_2205;
  reg  T_2207;
  reg [31:0] GEN_110;
  wire  T_2209;
  wire  T_2210;
  wire [1:0] T_2212;
  wire  T_2213;
  wire  GEN_54;
  wire  T_2215;
  wire  T_2216;
  wire [1:0] T_2218;
  wire  T_2219;
  wire  GEN_55;
  wire  T_2221;
  wire  T_2223;
  wire  T_2224;
  wire [25:0] GEN_56;
  wire [7:0] GEN_57;
  wire [3:0] GEN_58;
  wire  T_2231;
  wire  T_2233;
  wire  T_2234;
  wire  T_2236;
  wire  T_2237;
  wire  T_2239;
  wire  T_2240;
  wire  T_2241;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  wire  T_2251;
  wire [7:0] T_2252;
  wire  T_2253;
  wire  T_2254;
  wire  T_2255;
  wire  T_2256;
  wire  T_2257;
  wire  T_2263;
  wire  T_2264;
  wire  T_2266;
  wire  T_2267;
  wire  T_2271;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2286;
  wire  T_2288;
  wire  T_2289;
  wire [2:0] GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  T_2303;
  wire [7:0] T_2307;
  wire [7:0] T_2308;
  wire [7:0] T_2310;
  wire [7:0] T_2311;
  wire [7:0] T_2312;
  wire [7:0] T_2314;
  wire [2:0] GEN_62;
  wire  GEN_63;
  wire  GEN_64;
  wire [7:0] GEN_65;
  wire  T_2316;
  wire [7:0] T_2333;
  wire [7:0] GEN_66;
  wire [2:0] GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire [7:0] GEN_70;
  wire  T_2334;
  wire  T_2335;
  wire  T_2337;
  wire  T_2338;
  wire  T_2339;
  wire  T_2340;
  wire  T_2341;
  wire  T_2343;
  wire  T_2344;
  wire  T_2346;
  wire  T_2347;
  wire [2:0] T_2379_addr_beat;
  wire [25:0] T_2379_addr_block;
  wire  T_2379_client_xact_id;
  wire  T_2379_voluntary;
  wire [2:0] T_2379_r_type;
  wire [63:0] T_2379_data;
  wire  T_2379_client_id;
  wire [2:0] T_2440_addr_beat;
  wire  T_2440_client_xact_id;
  wire [1:0] T_2440_manager_xact_id;
  wire  T_2440_is_builtin_type;
  wire [3:0] T_2440_g_type;
  wire [63:0] T_2440_data;
  wire  T_2440_client_id;
  wire [7:0] GEN_0;
  wire [7:0] GEN_71;
  wire [7:0] GEN_72;
  wire [7:0] GEN_73;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire  T_2521;
  wire [7:0] GEN_1;
  wire  T_2522;
  wire [7:0] GEN_2;
  wire  T_2523;
  wire [7:0] GEN_3;
  wire  T_2524;
  wire [7:0] GEN_4;
  wire  T_2525;
  wire [7:0] GEN_5;
  wire  T_2526;
  wire [7:0] GEN_6;
  wire  T_2527;
  wire [7:0] GEN_7;
  wire  T_2528;
  wire [7:0] T_2532;
  wire [7:0] T_2536;
  wire [7:0] T_2540;
  wire [7:0] T_2544;
  wire [7:0] T_2548;
  wire [7:0] T_2552;
  wire [7:0] T_2556;
  wire [7:0] T_2560;
  wire [15:0] T_2561;
  wire [15:0] T_2562;
  wire [31:0] T_2563;
  wire [15:0] T_2564;
  wire [15:0] T_2565;
  wire [31:0] T_2566;
  wire [63:0] T_2567;
  wire [63:0] T_2568;
  wire [63:0] T_2569;
  wire [63:0] GEN_8;
  wire [63:0] GEN_127;
  wire [63:0] GEN_128;
  wire [63:0] GEN_129;
  wire [63:0] GEN_130;
  wire [63:0] GEN_131;
  wire [63:0] GEN_132;
  wire [63:0] GEN_133;
  wire [63:0] T_2570;
  wire [63:0] T_2571;
  wire [63:0] GEN_9;
  wire [63:0] GEN_134;
  wire [63:0] GEN_135;
  wire [63:0] GEN_136;
  wire [63:0] GEN_137;
  wire [63:0] GEN_138;
  wire [63:0] GEN_139;
  wire [63:0] GEN_140;
  wire [63:0] GEN_141;
  wire [7:0] GEN_10;
  wire [7:0] GEN_142;
  wire [7:0] GEN_143;
  wire [7:0] GEN_144;
  wire [7:0] GEN_145;
  wire [7:0] GEN_146;
  wire [7:0] GEN_147;
  wire [7:0] GEN_148;
  wire [7:0] GEN_149;
  wire [63:0] GEN_160;
  wire [63:0] GEN_161;
  wire [63:0] GEN_162;
  wire [63:0] GEN_163;
  wire [63:0] GEN_164;
  wire [63:0] GEN_165;
  wire [63:0] GEN_166;
  wire [63:0] GEN_167;
  wire [7:0] GEN_169;
  wire [7:0] GEN_170;
  wire [7:0] GEN_171;
  wire [7:0] GEN_172;
  wire [7:0] GEN_173;
  wire [7:0] GEN_174;
  wire [7:0] GEN_175;
  wire [7:0] GEN_176;
  wire [1:0] T_2604_state;
  wire  T_2631;
  wire [7:0] T_2647;
  wire [7:0] T_2648;
  wire  T_2651;
  wire  T_2652;
  wire  T_2653;
  wire  T_2654;
  wire  T_2655;
  wire  T_2656;
  wire [7:0] T_2660;
  wire [7:0] T_2661;
  wire [7:0] T_2663;
  wire [7:0] T_2664;
  wire [7:0] T_2665;
  wire [7:0] T_2666;
  wire [7:0] GEN_177;
  wire  T_2677;
  wire  T_2679;
  wire  T_2680;
  wire  GEN_179;
  wire  T_2692;
  wire  T_2693;
  wire  GEN_180;
  wire  GEN_181;
  wire  GEN_182;
  wire  T_2702;
  wire  T_2710;
  reg [2:0] T_2712;
  reg [31:0] GEN_111;
  wire  T_2714;
  wire [3:0] T_2716;
  wire [2:0] T_2717;
  wire [2:0] GEN_183;
  wire  T_2718;
  wire [2:0] T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [2:0] T_2733_0;
  wire [3:0] GEN_413;
  wire  T_2735;
  wire  T_2737;
  wire  T_2739;
  reg [2:0] T_2741;
  reg [31:0] GEN_112;
  wire  T_2743;
  wire [3:0] T_2745;
  wire [2:0] T_2746;
  wire [2:0] GEN_184;
  wire  T_2747;
  wire [2:0] T_2748;
  wire  T_2749;
  reg  T_2751;
  reg [31:0] GEN_113;
  wire  T_2753;
  wire  T_2754;
  wire [1:0] T_2756;
  wire  T_2757;
  wire  GEN_185;
  wire  T_2759;
  wire  T_2760;
  wire [1:0] T_2762;
  wire  T_2763;
  wire  GEN_186;
  wire  T_2765;
  wire [7:0] T_2774;
  wire  T_2775;
  wire  T_2776;
  wire  T_2777;
  wire  T_2791;
  wire [2:0] T_2792;
  wire [2:0] T_2828_addr_beat;
  wire [25:0] T_2828_addr_block;
  wire [1:0] T_2828_client_xact_id;
  wire  T_2828_voluntary;
  wire [2:0] T_2828_r_type;
  wire [63:0] T_2828_data;
  wire [63:0] GEN_11;
  wire [63:0] GEN_187;
  wire [63:0] GEN_188;
  wire [63:0] GEN_189;
  wire [63:0] GEN_190;
  wire [63:0] GEN_191;
  wire [63:0] GEN_192;
  wire [63:0] GEN_193;
  wire  T_2857;
  wire  T_2860;
  wire [2:0] T_2871_0;
  wire  T_2873;
  wire  T_2874;
  wire  T_2875;
  reg [2:0] T_2877;
  reg [31:0] GEN_114;
  wire  T_2879;
  wire [3:0] T_2881;
  wire [2:0] T_2882;
  wire [2:0] GEN_195;
  wire  T_2883;
  wire [2:0] T_2884;
  wire  T_2885;
  wire  T_2891;
  wire  T_2892;
  wire [2:0] T_2900_0;
  wire [3:0] GEN_414;
  wire  T_2902;
  wire  T_2904;
  wire  T_2906;
  reg [2:0] T_2908;
  reg [31:0] GEN_115;
  wire  T_2910;
  wire [3:0] T_2912;
  wire [2:0] T_2913;
  wire [2:0] GEN_196;
  wire  T_2914;
  wire [2:0] T_2915;
  wire  T_2916;
  reg  T_2918;
  reg [31:0] GEN_116;
  wire  T_2920;
  wire  T_2921;
  wire [1:0] T_2923;
  wire  T_2924;
  wire  GEN_197;
  wire  T_2926;
  wire  T_2927;
  wire [1:0] T_2929;
  wire  T_2930;
  wire  GEN_198;
  wire  T_2932;
  wire  T_2933;
  wire [7:0] T_2937;
  wire  T_2938;
  wire  T_2940;
  wire [2:0] T_2949_0;
  wire [2:0] T_2949_1;
  wire [2:0] T_2949_2;
  wire  T_2967;
  wire  T_2968;
  wire  T_2971;
  wire  T_2972;
  wire  T_2973;
  wire  T_2974;
  wire  T_2975;
  wire  T_2976;
  wire  T_2977;
  wire  T_2978;
  wire  T_2979;
  wire  T_2980;
  wire  T_2981;
  wire [5:0] T_2984;
  wire [25:0] T_3015_addr_block;
  wire [1:0] T_3015_client_xact_id;
  wire [2:0] T_3015_addr_beat;
  wire  T_3015_is_builtin_type;
  wire [2:0] T_3015_a_type;
  wire [10:0] T_3015_union;
  wire [63:0] T_3015_data;
  wire [7:0] GEN_12;
  wire [7:0] GEN_199;
  wire [7:0] GEN_200;
  wire [7:0] GEN_201;
  wire [7:0] GEN_202;
  wire [7:0] GEN_203;
  wire [7:0] GEN_204;
  wire [7:0] GEN_205;
  wire [5:0] T_3080;
  wire [4:0] T_3081;
  wire [10:0] T_3082;
  wire [6:0] T_3084;
  wire [7:0] T_3085;
  wire [8:0] T_3087;
  wire [5:0] T_3099;
  wire [5:0] T_3101;
  wire [10:0] T_3103;
  wire [10:0] T_3105;
  wire [10:0] T_3107;
  wire [10:0] T_3109;
  wire [10:0] T_3111;
  wire [25:0] T_3140_addr_block;
  wire [1:0] T_3140_client_xact_id;
  wire [2:0] T_3140_addr_beat;
  wire  T_3140_is_builtin_type;
  wire [2:0] T_3140_a_type;
  wire [10:0] T_3140_union;
  wire [63:0] T_3140_data;
  wire [63:0] GEN_13;
  wire [63:0] GEN_206;
  wire [63:0] GEN_207;
  wire [63:0] GEN_208;
  wire [63:0] GEN_209;
  wire [63:0] GEN_210;
  wire [63:0] GEN_211;
  wire [63:0] GEN_212;
  wire [25:0] T_3168_addr_block;
  wire [1:0] T_3168_client_xact_id;
  wire [2:0] T_3168_addr_beat;
  wire  T_3168_is_builtin_type;
  wire [2:0] T_3168_a_type;
  wire [10:0] T_3168_union;
  wire [63:0] T_3168_data;
  wire  T_3197;
  wire [3:0] GEN_213;
  wire  GEN_214;
  wire [2:0] T_3207_0;
  wire [2:0] T_3207_1;
  wire [3:0] GEN_415;
  wire  T_3209;
  wire [3:0] GEN_416;
  wire  T_3210;
  wire  T_3211;
  wire  T_3213;
  wire  T_3214;
  wire [7:0] GEN_14;
  wire [7:0] GEN_215;
  wire [7:0] GEN_216;
  wire [7:0] GEN_217;
  wire [7:0] GEN_218;
  wire [7:0] GEN_219;
  wire [7:0] GEN_220;
  wire [7:0] GEN_221;
  wire  T_3215;
  wire [7:0] GEN_15;
  wire  T_3216;
  wire [7:0] GEN_16;
  wire  T_3217;
  wire [7:0] GEN_17;
  wire  T_3218;
  wire [7:0] GEN_18;
  wire  T_3219;
  wire [7:0] GEN_19;
  wire  T_3220;
  wire [7:0] GEN_20;
  wire  T_3221;
  wire [7:0] GEN_21;
  wire  T_3222;
  wire [7:0] T_3226;
  wire [7:0] T_3230;
  wire [7:0] T_3234;
  wire [7:0] T_3238;
  wire [7:0] T_3242;
  wire [7:0] T_3246;
  wire [7:0] T_3250;
  wire [7:0] T_3254;
  wire [15:0] T_3255;
  wire [15:0] T_3256;
  wire [31:0] T_3257;
  wire [15:0] T_3258;
  wire [15:0] T_3259;
  wire [31:0] T_3260;
  wire [63:0] T_3261;
  wire [63:0] T_3262;
  wire [63:0] T_3263;
  wire [63:0] GEN_22;
  wire [63:0] GEN_271;
  wire [63:0] GEN_272;
  wire [63:0] GEN_273;
  wire [63:0] GEN_274;
  wire [63:0] GEN_275;
  wire [63:0] GEN_276;
  wire [63:0] GEN_277;
  wire [63:0] T_3264;
  wire [63:0] T_3265;
  wire [63:0] GEN_23;
  wire [63:0] GEN_278;
  wire [63:0] GEN_279;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [7:0] GEN_24;
  wire [7:0] GEN_286;
  wire [7:0] GEN_287;
  wire [7:0] GEN_288;
  wire [7:0] GEN_289;
  wire [7:0] GEN_290;
  wire [7:0] GEN_291;
  wire [7:0] GEN_292;
  wire [7:0] GEN_293;
  wire [63:0] GEN_304;
  wire [63:0] GEN_305;
  wire [63:0] GEN_306;
  wire [63:0] GEN_307;
  wire [63:0] GEN_308;
  wire [63:0] GEN_309;
  wire [63:0] GEN_310;
  wire [63:0] GEN_311;
  wire [7:0] GEN_313;
  wire [7:0] GEN_314;
  wire [7:0] GEN_315;
  wire [7:0] GEN_316;
  wire [7:0] GEN_317;
  wire [7:0] GEN_318;
  wire [7:0] GEN_319;
  wire [7:0] GEN_320;
  wire  T_3268;
  wire  T_3269;
  wire  T_3281;
  wire  T_3283;
  wire [2:0] T_3291_0;
  wire [3:0] GEN_417;
  wire  T_3293;
  wire  T_3295;
  wire  T_3297;
  reg [2:0] T_3299;
  reg [31:0] GEN_117;
  wire  T_3301;
  wire [3:0] T_3303;
  wire [2:0] T_3304;
  wire [2:0] GEN_321;
  wire  T_3305;
  wire [2:0] T_3306;
  wire  T_3307;
  wire  T_3308;
  reg [2:0] T_3314;
  reg [31:0] GEN_118;
  reg  T_3324;
  reg [31:0] GEN_119;
  wire  T_3326;
  wire  T_3327;
  wire [1:0] T_3329;
  wire  T_3330;
  wire  GEN_323;
  wire  T_3332;
  wire  T_3333;
  wire [1:0] T_3335;
  wire  T_3336;
  wire  GEN_324;
  wire  T_3338;
  wire  T_3343;
  wire [7:0] T_3360;
  wire [2:0] T_3370_0;
  wire [2:0] T_3370_1;
  wire [3:0] GEN_418;
  wire  T_3372;
  wire [3:0] GEN_419;
  wire  T_3373;
  wire  T_3374;
  wire  T_3376;
  wire  T_3377;
  wire [7:0] T_3382;
  wire [7:0] T_3384;
  wire [7:0] T_3385;
  wire [7:0] T_3386;
  wire [7:0] GEN_327;
  wire  T_3389;
  wire  T_3390;
  wire  T_3393;
  wire  T_3395;
  wire  T_3412;
  wire [2:0] T_3413;
  wire  T_3414;
  wire [2:0] T_3415;
  wire  T_3416;
  wire [2:0] T_3417;
  wire  T_3418;
  wire [2:0] T_3419;
  wire  T_3420;
  wire [2:0] T_3421;
  wire  T_3422;
  wire [2:0] T_3423;
  wire  T_3424;
  wire [2:0] T_3425;
  wire [2:0] T_3426;
  wire [2:0] T_3455_addr_beat;
  wire  T_3455_client_xact_id;
  wire [1:0] T_3455_manager_xact_id;
  wire  T_3455_is_builtin_type;
  wire [3:0] T_3455_g_type;
  wire [63:0] T_3455_data;
  wire  T_3455_client_id;
  wire [63:0] GEN_25;
  wire [63:0] GEN_328;
  wire [63:0] GEN_329;
  wire [63:0] GEN_330;
  wire [63:0] GEN_331;
  wire [63:0] GEN_332;
  wire [63:0] GEN_333;
  wire [63:0] GEN_334;
  wire [2:0] T_3491_0;
  wire [3:0] GEN_420;
  wire  T_3493;
  wire  T_3495;
  wire  T_3497;
  reg [2:0] T_3499;
  reg [31:0] GEN_120;
  wire  T_3501;
  wire [3:0] T_3503;
  wire [2:0] T_3504;
  wire [2:0] GEN_335;
  wire  T_3505;
  wire [2:0] T_3506;
  wire  T_3507;
  wire  T_3512;
  wire  T_3514;
  wire [2:0] T_3522_0;
  wire [2:0] T_3522_1;
  wire [3:0] GEN_421;
  wire  T_3524;
  wire [3:0] GEN_422;
  wire  T_3525;
  wire  T_3526;
  wire  T_3528;
  wire [7:0] T_3529;
  wire  T_3530;
  wire  T_3532;
  wire  T_3533;
  wire  GEN_338;
  wire  GEN_339;
  wire [2:0] GEN_340;
  wire  GEN_341;
  wire [1:0] GEN_342;
  wire  GEN_343;
  wire [3:0] GEN_344;
  wire [63:0] GEN_345;
  wire  GEN_346;
  wire  GEN_349;
  wire  T_3540;
  wire [1:0] GEN_350;
  wire  T_3551;
  wire  T_3552;
  wire [2:0] T_3562_0;
  wire [2:0] T_3562_1;
  wire [2:0] T_3562_2;
  wire  T_3564;
  wire  T_3565;
  wire  T_3566;
  wire  T_3567;
  wire  T_3568;
  wire  T_3569;
  wire  T_3570;
  wire  T_3571;
  wire  T_3573;
  wire  T_3574;
  wire  T_3603;
  wire [7:0] T_3604;
  wire [7:0] T_3606;
  wire [7:0] T_3607;
  wire  T_3608;
  wire  T_3609;
  wire  T_3610;
  wire  T_3611;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3615;
  wire [7:0] T_3619;
  wire [7:0] T_3623;
  wire [7:0] T_3627;
  wire [7:0] T_3631;
  wire [7:0] T_3635;
  wire [7:0] T_3639;
  wire [7:0] T_3643;
  wire [7:0] T_3647;
  wire [15:0] T_3648;
  wire [15:0] T_3649;
  wire [31:0] T_3650;
  wire [15:0] T_3651;
  wire [15:0] T_3652;
  wire [31:0] T_3653;
  wire [63:0] T_3654;
  wire [63:0] T_3655;
  wire [63:0] GEN_26;
  wire [63:0] GEN_351;
  wire [63:0] GEN_352;
  wire [63:0] GEN_353;
  wire [63:0] GEN_354;
  wire [63:0] GEN_355;
  wire [63:0] GEN_356;
  wire [63:0] GEN_357;
  wire [63:0] T_3656;
  wire [63:0] T_3657;
  wire [63:0] T_3658;
  wire [63:0] GEN_27;
  wire [63:0] GEN_358;
  wire [63:0] GEN_359;
  wire [63:0] GEN_360;
  wire [63:0] GEN_361;
  wire [63:0] GEN_362;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [7:0] GEN_28;
  wire [7:0] GEN_366;
  wire [7:0] GEN_367;
  wire [7:0] GEN_368;
  wire [7:0] GEN_369;
  wire [7:0] GEN_370;
  wire [7:0] GEN_371;
  wire [7:0] GEN_372;
  wire [7:0] T_3695;
  wire [7:0] GEN_29;
  wire [7:0] GEN_373;
  wire [7:0] GEN_374;
  wire [7:0] GEN_375;
  wire [7:0] GEN_376;
  wire [7:0] GEN_377;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [63:0] GEN_383;
  wire [63:0] GEN_384;
  wire [63:0] GEN_385;
  wire [63:0] GEN_386;
  wire [63:0] GEN_387;
  wire [63:0] GEN_388;
  wire [63:0] GEN_389;
  wire [63:0] GEN_390;
  wire [7:0] GEN_393;
  wire [7:0] GEN_394;
  wire [7:0] GEN_395;
  wire [7:0] GEN_396;
  wire [7:0] GEN_397;
  wire [7:0] GEN_398;
  wire [7:0] GEN_399;
  wire [7:0] GEN_400;
  wire  T_3698;
  wire  T_3699;
  wire  T_3700;
  wire  T_3701;
  wire  T_3702;
  wire  T_3703;
  wire  T_3704;
  wire  T_3706;
  wire  T_3708;
  wire [3:0] GEN_401;
  wire [7:0] GEN_402;
  wire [7:0] GEN_403;
  wire [7:0] GEN_404;
  wire [7:0] GEN_405;
  wire [7:0] GEN_406;
  wire [7:0] GEN_407;
  wire [7:0] GEN_408;
  wire [7:0] GEN_409;
  wire  GEN_30;
  reg [31:0] GEN_121;
  wire  GEN_31;
  reg [31:0] GEN_122;
  Queue_8 ignt_q (
    .clk(ignt_q_clk),
    .reset(ignt_q_reset),
    .io_enq_ready(ignt_q_io_enq_ready),
    .io_enq_valid(ignt_q_io_enq_valid),
    .io_enq_bits_client_xact_id(ignt_q_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(ignt_q_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(ignt_q_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(ignt_q_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(ignt_q_io_enq_bits_a_type),
    .io_deq_ready(ignt_q_io_deq_ready),
    .io_deq_valid(ignt_q_io_deq_valid),
    .io_deq_bits_client_xact_id(ignt_q_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(ignt_q_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(ignt_q_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(ignt_q_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(ignt_q_io_deq_bits_a_type),
    .io_count(ignt_q_io_count)
  );
  assign io_inner_acquire_ready = T_1981;
  assign io_inner_grant_valid = GEN_349;
  assign io_inner_grant_bits_addr_beat = GEN_340;
  assign io_inner_grant_bits_client_xact_id = GEN_341;
  assign io_inner_grant_bits_manager_xact_id = GEN_342;
  assign io_inner_grant_bits_is_builtin_type = GEN_343;
  assign io_inner_grant_bits_g_type = GEN_344;
  assign io_inner_grant_bits_data = GEN_345;
  assign io_inner_grant_bits_client_id = GEN_346;
  assign io_inner_finish_ready = T_2337;
  assign io_inner_probe_valid = T_2083;
  assign io_inner_probe_bits_addr_block = T_2030_addr_block;
  assign io_inner_probe_bits_p_type = T_2030_p_type;
  assign io_inner_probe_bits_client_id = T_2030_client_id;
  assign io_inner_release_ready = T_2274;
  assign io_outer_acquire_valid = T_2968;
  assign io_outer_acquire_bits_addr_block = T_3168_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3168_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3168_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3168_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3168_a_type;
  assign io_outer_acquire_bits_union = T_3168_union;
  assign io_outer_acquire_bits_data = T_3168_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2777;
  assign io_outer_release_bits_addr_beat = T_2828_addr_beat;
  assign io_outer_release_bits_addr_block = T_2828_addr_block;
  assign io_outer_release_bits_client_xact_id = T_2828_client_xact_id;
  assign io_outer_release_bits_voluntary = T_2828_voluntary;
  assign io_outer_release_bits_r_type = T_2828_r_type;
  assign io_outer_release_bits_data = T_2828_data;
  assign io_outer_grant_ready = GEN_214;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_30;
  assign io_outer_finish_bits_manager_id = GEN_31;
  assign io_alloc_iacq_matches = T_1749;
  assign io_alloc_iacq_can = T_1611;
  assign io_alloc_irel_matches = T_1752;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1755;
  assign io_alloc_oprb_can = 1'h0;
  assign io_alloc_idle = T_1611;
  assign io_alloc_addr_block = xact_addr_block;
  assign all_pending_done = T_3706;
  assign xact_addr_beat = xact_iacq_addr_beat;
  assign xact_iacq_client_xact_id = T_1823_client_xact_id;
  assign xact_iacq_addr_beat = T_1823_addr_beat;
  assign xact_iacq_client_id = T_1823_client_id;
  assign xact_iacq_is_builtin_type = T_1823_is_builtin_type;
  assign xact_iacq_a_type = T_1823_a_type;
  assign vol_ignt_counter_pending = T_2221;
  assign vol_ignt_counter_up_idx = T_2173;
  assign vol_ignt_counter_up_done = T_2174;
  assign vol_ignt_counter_down_idx = T_2204;
  assign vol_ignt_counter_down_done = T_2205;
  assign scoreboard_6 = T_1850;
  assign ignt_data_idx = T_3506;
  assign ignt_data_done = T_3507;
  assign ifin_counter_pending = T_3338;
  assign ifin_counter_up_idx = T_3306;
  assign ifin_counter_up_done = T_3307;
  assign ifin_counter_down_idx = 3'h0;
  assign ifin_counter_down_done = T_3308;
  assign ognt_counter_pending = T_2932;
  assign ognt_counter_up_idx = T_2884;
  assign ognt_counter_up_done = T_2885;
  assign ognt_counter_down_idx = T_2915;
  assign ognt_counter_down_done = T_2916;
  assign vol_ognt_counter_pending = T_2765;
  assign vol_ognt_counter_up_idx = T_2719;
  assign vol_ognt_counter_up_done = T_2720;
  assign vol_ognt_counter_down_idx = T_2748;
  assign vol_ognt_counter_down_done = T_2749;
  assign T_170 = pending_orel_data != 8'h0;
  assign T_171 = pending_orel_send | T_170;
  assign scoreboard_3 = T_171 | vol_ognt_counter_pending;
  assign T_195_sharers = 1'h0;
  assign T_241_state = 2'h0;
  assign coh_inner_sharers = T_195_sharers;
  assign coh_outer_state = T_241_state;
  assign T_1611 = state == 4'h0;
  assign T_1612 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1613 = T_1611 & T_1612;
  assign T_1614 = T_1613 & io_alloc_iacq_should;
  assign T_1623_0 = 3'h3;
  assign T_1625 = io_inner_acquire_bits_a_type == T_1623_0;
  assign T_1626 = io_inner_acquire_bits_is_builtin_type & T_1625;
  assign T_1627 = T_1614 & T_1626;
  assign T_1636_0 = 3'h3;
  assign T_1638 = io_inner_acquire_bits_a_type == T_1636_0;
  assign T_1639 = io_inner_acquire_bits_is_builtin_type & T_1638;
  assign T_1641 = T_1639 == 1'h0;
  assign T_1643 = io_inner_acquire_bits_addr_beat == 3'h0;
  assign T_1644 = T_1641 | T_1643;
  assign T_1646 = T_1644 == 1'h0;
  assign T_1647 = T_1627 & T_1646;
  assign T_1649 = T_1647 == 1'h0;
  assign T_1650 = T_1649 | reset;
  assign T_1652 = T_1650 == 1'h0;
  assign T_1653 = state != 4'h0;
  assign T_1654 = T_1653 & scoreboard_6;
  assign T_1656 = xact_iacq_a_type == 3'h5;
  assign T_1658 = xact_iacq_a_type == 3'h6;
  assign T_1659 = T_1656 | T_1658;
  assign T_1660 = xact_iacq_is_builtin_type & T_1659;
  assign T_1661 = T_1654 & T_1660;
  assign T_1663 = T_1661 == 1'h0;
  assign T_1664 = T_1663 | reset;
  assign T_1666 = T_1664 == 1'h0;
  assign T_1670 = xact_iacq_a_type == 3'h4;
  assign T_1671 = xact_iacq_is_builtin_type & T_1670;
  assign T_1672 = T_1654 & T_1671;
  assign T_1674 = T_1672 == 1'h0;
  assign T_1675 = T_1674 | reset;
  assign T_1677 = T_1675 == 1'h0;
  assign T_1691_0 = 64'h0;
  assign T_1691_1 = 64'h0;
  assign T_1691_2 = 64'h0;
  assign T_1691_3 = 64'h0;
  assign T_1691_4 = 64'h0;
  assign T_1691_5 = 64'h0;
  assign T_1691_6 = 64'h0;
  assign T_1691_7 = 64'h0;
  assign T_1709_0 = 8'h0;
  assign T_1709_1 = 8'h0;
  assign T_1709_2 = 8'h0;
  assign T_1709_3 = 8'h0;
  assign T_1709_4 = 8'h0;
  assign T_1709_5 = 8'h0;
  assign T_1709_6 = 8'h0;
  assign T_1709_7 = 8'h0;
  assign T_1714 = ~ wmask_buffer_0;
  assign T_1716 = T_1714 == 8'h0;
  assign T_1717 = ~ wmask_buffer_1;
  assign T_1719 = T_1717 == 8'h0;
  assign T_1720 = ~ wmask_buffer_2;
  assign T_1722 = T_1720 == 8'h0;
  assign T_1723 = ~ wmask_buffer_3;
  assign T_1725 = T_1723 == 8'h0;
  assign T_1726 = ~ wmask_buffer_4;
  assign T_1728 = T_1726 == 8'h0;
  assign T_1729 = ~ wmask_buffer_5;
  assign T_1731 = T_1729 == 8'h0;
  assign T_1732 = ~ wmask_buffer_6;
  assign T_1734 = T_1732 == 8'h0;
  assign T_1735 = ~ wmask_buffer_7;
  assign T_1737 = T_1735 == 8'h0;
  assign data_valid_0 = T_1716;
  assign data_valid_1 = T_1719;
  assign data_valid_2 = T_1722;
  assign data_valid_3 = T_1725;
  assign data_valid_4 = T_1728;
  assign data_valid_5 = T_1731;
  assign data_valid_6 = T_1734;
  assign data_valid_7 = T_1737;
  assign T_1748 = io_inner_acquire_bits_addr_block == xact_addr_block;
  assign T_1749 = T_1653 & T_1748;
  assign T_1751 = io_inner_release_bits_addr_block == xact_addr_block;
  assign T_1752 = T_1653 & T_1751;
  assign T_1754 = io_outer_probe_bits_addr_block == xact_addr_block;
  assign T_1755 = T_1653 & T_1754;
  assign T_1764 = xact_iacq_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1765 = xact_iacq_client_id == io_inner_acquire_bits_client_id;
  assign T_1766 = T_1764 & T_1765;
  assign T_1767 = T_1766 & scoreboard_6;
  assign T_1768 = xact_iacq_addr_beat == io_inner_acquire_bits_addr_beat;
  assign T_1769 = T_1767 & T_1768;
  assign ignt_q_clk = clk;
  assign ignt_q_reset = reset;
  assign ignt_q_io_enq_valid = T_1822;
  assign ignt_q_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign ignt_q_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign ignt_q_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign ignt_q_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign ignt_q_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign ignt_q_io_deq_ready = GEN_339;
  assign T_1797 = T_1611 & io_alloc_iacq_should;
  assign T_1798 = T_1797 & io_inner_acquire_valid;
  assign T_1800 = T_1769 == 1'h0;
  assign T_1801 = T_1800 & scoreboard_6;
  assign T_1803 = T_1801 & T_1612;
  assign T_1812_0 = 3'h3;
  assign T_1814 = io_inner_acquire_bits_a_type == T_1812_0;
  assign T_1815 = io_inner_acquire_bits_is_builtin_type & T_1814;
  assign T_1817 = T_1815 == 1'h0;
  assign T_1820 = T_1817 | T_1643;
  assign T_1821 = T_1803 & T_1820;
  assign T_1822 = T_1798 | T_1821;
  assign T_1823_client_xact_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_xact_id : ignt_q_io_enq_bits_client_xact_id;
  assign T_1823_addr_beat = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_addr_beat : ignt_q_io_enq_bits_addr_beat;
  assign T_1823_client_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_id : ignt_q_io_enq_bits_client_id;
  assign T_1823_is_builtin_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_is_builtin_type : ignt_q_io_enq_bits_is_builtin_type;
  assign T_1823_a_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_a_type : ignt_q_io_enq_bits_a_type;
  assign T_1850 = ignt_q_io_count > 2'h0;
  assign T_1852 = T_1653 | io_alloc_iacq_should;
  assign T_1862_0 = 3'h2;
  assign T_1862_1 = 3'h3;
  assign T_1862_2 = 3'h4;
  assign T_1864 = io_inner_acquire_bits_a_type == T_1862_0;
  assign T_1865 = io_inner_acquire_bits_a_type == T_1862_1;
  assign T_1866 = io_inner_acquire_bits_a_type == T_1862_2;
  assign T_1867 = T_1864 | T_1865;
  assign T_1868 = T_1867 | T_1866;
  assign T_1869 = io_inner_acquire_bits_is_builtin_type & T_1868;
  assign T_1870 = T_1612 & T_1869;
  assign T_1874 = T_1870 ? 8'hff : 8'h0;
  assign T_1875 = ~ T_1874;
  assign T_1877 = 8'h1 << io_inner_acquire_bits_addr_beat;
  assign T_1878 = ~ T_1877;
  assign T_1879 = T_1875 | T_1878;
  assign T_1880 = pending_put_data & T_1879;
  assign T_1890_0 = 3'h3;
  assign T_1892 = io_inner_acquire_bits_a_type == T_1890_0;
  assign T_1893 = io_inner_acquire_bits_is_builtin_type & T_1892;
  assign T_1894 = T_1612 & T_1893;
  assign T_1897 = T_1894 & T_1643;
  assign T_1906 = T_1897 ? 8'hfe : 8'h0;
  assign T_1907 = T_1880 | T_1906;
  assign GEN_34 = T_1852 ? T_1907 : pending_put_data;
  assign T_1915 = 4'h8 * 4'h0;
  assign T_1917 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1918 = io_inner_acquire_bits_is_builtin_type & T_1917;
  assign T_1920 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1921 = io_inner_acquire_bits_is_builtin_type & T_1920;
  assign T_1922 = T_1918 | T_1921;
  assign T_1923 = io_inner_acquire_bits_union[5:1];
  assign T_1924 = T_1922 ? 5'h1 : T_1923;
  assign T_1925 = io_inner_acquire_bits_union[10:8];
  assign T_1926 = io_inner_acquire_bits_union[7:6];
  assign T_1939_0 = 3'h2;
  assign T_1939_1 = 3'h3;
  assign T_1939_2 = 3'h4;
  assign T_1941 = io_inner_acquire_bits_a_type == T_1939_0;
  assign T_1942 = io_inner_acquire_bits_a_type == T_1939_1;
  assign T_1943 = io_inner_acquire_bits_a_type == T_1939_2;
  assign T_1944 = T_1941 | T_1942;
  assign T_1945 = T_1944 | T_1943;
  assign T_1946 = io_inner_acquire_bits_is_builtin_type & T_1945;
  assign T_1947 = T_1612 & T_1946;
  assign T_1951 = T_1947 ? 8'hff : 8'h0;
  assign T_1952 = ~ T_1951;
  assign T_1956 = T_1952 | T_1878;
  assign T_1958 = T_1921 ? T_1956 : 8'h0;
  assign GEN_35 = T_1798 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_36 = T_1798 ? 1'h0 : xact_allocate;
  assign GEN_37 = T_1798 ? T_1915 : xact_amo_shift_bytes;
  assign GEN_38 = T_1798 ? T_1924 : xact_op_code;
  assign GEN_39 = T_1798 ? T_1925 : xact_addr_byte;
  assign GEN_40 = T_1798 ? T_1926 : xact_op_size;
  assign GEN_44 = T_1798 ? T_1958 : GEN_34;
  assign GEN_45 = T_1798 ? 8'h0 : pending_ignt_data;
  assign GEN_46 = T_1798 ? 4'h5 : state;
  assign scoreboard_0 = pending_put_data != 8'h0;
  assign T_1976_0 = 3'h3;
  assign T_1978 = io_inner_acquire_bits_a_type == T_1976_0;
  assign T_1979 = io_inner_acquire_bits_is_builtin_type & T_1978;
  assign T_1980 = T_1767 & T_1979;
  assign T_1981 = T_1611 | T_1980;
  assign T_1982 = ~ pending_ignt_data;
  assign skip_outer_acquire = T_1982 == 8'h0;
  assign T_1991 = 3'h4 == xact_iacq_a_type;
  assign T_1992 = T_1991 ? 2'h0 : 2'h2;
  assign T_1993 = 3'h6 == xact_iacq_a_type;
  assign T_1994 = T_1993 ? 2'h0 : T_1992;
  assign T_1995 = 3'h5 == xact_iacq_a_type;
  assign T_1996 = T_1995 ? 2'h2 : T_1994;
  assign T_1997 = 3'h2 == xact_iacq_a_type;
  assign T_1998 = T_1997 ? 2'h0 : T_1996;
  assign T_1999 = 3'h0 == xact_iacq_a_type;
  assign T_2000 = T_1999 ? 2'h2 : T_1998;
  assign T_2001 = 3'h3 == xact_iacq_a_type;
  assign T_2002 = T_2001 ? 2'h0 : T_2000;
  assign T_2003 = 3'h1 == xact_iacq_a_type;
  assign T_2004 = T_2003 ? 2'h2 : T_2002;
  assign T_2005 = xact_iacq_is_builtin_type ? T_2004 : 2'h0;
  assign T_2030_addr_block = xact_addr_block;
  assign T_2030_p_type = T_2005;
  assign T_2030_client_id = 1'h0;
  assign T_2055 = skip_outer_acquire == 1'h0;
  assign T_2056 = T_2055 ? 4'h6 : 4'h7;
  assign T_2065_pending = T_2139;
  assign T_2065_up_idx = 3'h0;
  assign T_2065_up_done = T_2073;
  assign T_2065_down_idx = T_2122;
  assign T_2065_down_done = T_2123;
  assign T_2073 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2074 = ~ T_2073;
  assign T_2076 = 2'h1 << io_inner_probe_bits_client_id;
  assign T_2077 = ~ T_2076;
  assign GEN_410 = {{1'd0}, T_2074};
  assign T_2078 = GEN_410 | T_2077;
  assign GEN_411 = {{1'd0}, pending_iprbs};
  assign T_2079 = GEN_411 & T_2078;
  assign T_2080 = state == 4'h5;
  assign T_2083 = T_2080 & pending_iprbs;
  assign T_2100 = io_inner_release_ready & io_inner_release_valid;
  assign T_2103 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2104 = T_1653 & T_2103;
  assign T_2105 = T_2100 & T_2104;
  assign T_2107 = io_inner_release_bits_r_type == 3'h0;
  assign T_2108 = io_inner_release_bits_r_type == 3'h1;
  assign T_2109 = io_inner_release_bits_r_type == 3'h2;
  assign T_2110 = T_2107 | T_2108;
  assign T_2111 = T_2110 | T_2109;
  assign T_2113 = T_2105 & T_2111;
  assign T_2117 = T_2115 == 3'h7;
  assign T_2119 = T_2115 + 3'h1;
  assign T_2120 = T_2119[2:0];
  assign GEN_48 = T_2113 ? T_2120 : T_2115;
  assign T_2121 = T_2113 & T_2117;
  assign T_2122 = T_2111 ? T_2115 : 3'h0;
  assign T_2123 = T_2111 ? T_2121 : T_2105;
  assign T_2127 = T_2123 == 1'h0;
  assign T_2128 = T_2073 & T_2127;
  assign T_2130 = T_2125 + 1'h1;
  assign T_2131 = T_2130[0:0];
  assign GEN_49 = T_2128 ? T_2131 : T_2125;
  assign T_2133 = T_2073 == 1'h0;
  assign T_2134 = T_2123 & T_2133;
  assign T_2136 = T_2125 - 1'h1;
  assign T_2137 = T_2136[0:0];
  assign GEN_50 = T_2134 ? T_2137 : GEN_49;
  assign T_2139 = T_2125 > 1'h0;
  assign T_2143 = pending_iprbs | T_2065_pending;
  assign T_2145 = T_2143 == 1'h0;
  assign T_2146 = T_2080 & T_2145;
  assign GEN_51 = T_2146 ? T_2056 : GEN_46;
  assign T_2150 = T_1611 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2151 = T_2150 & io_inner_release_bits_voluntary;
  assign T_2156 = T_2100 & T_2151;
  assign T_2164 = T_2156 & T_2111;
  assign T_2168 = T_2166 == 3'h7;
  assign T_2170 = T_2166 + 3'h1;
  assign T_2171 = T_2170[2:0];
  assign GEN_52 = T_2164 ? T_2171 : T_2166;
  assign T_2172 = T_2164 & T_2168;
  assign T_2173 = T_2111 ? T_2166 : 3'h0;
  assign T_2174 = T_2111 ? T_2172 : T_2156;
  assign T_2175 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_2178 = io_inner_grant_bits_g_type == 4'h0;
  assign T_2179 = io_inner_grant_bits_is_builtin_type & T_2178;
  assign T_2180 = T_1653 & T_2179;
  assign T_2181 = T_2175 & T_2180;
  assign T_2189_0 = 3'h5;
  assign GEN_412 = {{1'd0}, T_2189_0};
  assign T_2191 = io_inner_grant_bits_g_type == GEN_412;
  assign T_2193 = io_inner_grant_bits_is_builtin_type ? T_2191 : T_2178;
  assign T_2195 = T_2181 & T_2193;
  assign T_2199 = T_2197 == 3'h7;
  assign T_2201 = T_2197 + 3'h1;
  assign T_2202 = T_2201[2:0];
  assign GEN_53 = T_2195 ? T_2202 : T_2197;
  assign T_2203 = T_2195 & T_2199;
  assign T_2204 = T_2193 ? T_2197 : 3'h0;
  assign T_2205 = T_2193 ? T_2203 : T_2181;
  assign T_2209 = T_2205 == 1'h0;
  assign T_2210 = T_2174 & T_2209;
  assign T_2212 = T_2207 + 1'h1;
  assign T_2213 = T_2212[0:0];
  assign GEN_54 = T_2210 ? T_2213 : T_2207;
  assign T_2215 = T_2174 == 1'h0;
  assign T_2216 = T_2205 & T_2215;
  assign T_2218 = T_2207 - 1'h1;
  assign T_2219 = T_2218[0:0];
  assign GEN_55 = T_2216 ? T_2219 : GEN_54;
  assign T_2221 = T_2207 > 1'h0;
  assign T_2223 = T_1611 & io_alloc_irel_should;
  assign T_2224 = T_2223 & io_inner_release_valid;
  assign GEN_56 = T_2224 ? io_inner_release_bits_addr_block : GEN_35;
  assign GEN_57 = T_2224 ? 8'hff : pending_irel_data;
  assign GEN_58 = T_2224 ? 4'h7 : GEN_51;
  assign T_2231 = T_1751 & io_inner_release_bits_voluntary;
  assign T_2233 = state == 4'h8;
  assign T_2234 = T_1611 | T_2233;
  assign T_2236 = T_2234 == 1'h0;
  assign T_2237 = T_2231 & T_2236;
  assign T_2239 = all_pending_done == 1'h0;
  assign T_2240 = T_2237 & T_2239;
  assign T_2241 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2243 = T_2241 == 1'h0;
  assign T_2244 = T_2240 & T_2243;
  assign T_2247 = T_2175 == 1'h0;
  assign T_2248 = T_2244 & T_2247;
  assign T_2250 = vol_ignt_counter_pending == 1'h0;
  assign T_2251 = T_2248 & T_2250;
  assign T_2252 = pending_orel_data >> io_inner_release_bits_addr_beat;
  assign T_2253 = T_2252[0];
  assign T_2254 = sending_orel & T_2253;
  assign T_2255 = io_outer_release_ready & io_outer_release_valid;
  assign T_2256 = io_inner_release_bits_addr_beat == io_outer_release_bits_addr_beat;
  assign T_2257 = T_2255 & T_2256;
  assign T_2263 = T_2254 | T_2257;
  assign T_2264 = T_2111 & T_2263;
  assign T_2266 = T_2264 == 1'h0;
  assign T_2267 = T_2251 & T_2266;
  assign T_2271 = T_1751 & T_2103;
  assign T_2273 = T_2271 & T_2080;
  assign T_2274 = T_2267 | T_2273;
  assign T_2275 = T_2274 & io_inner_release_valid;
  assign T_2276 = T_2224 | T_2275;
  assign T_2277 = T_2276 & io_inner_release_ready;
  assign T_2286 = T_2111 == 1'h0;
  assign T_2288 = io_inner_release_bits_addr_beat == 3'h0;
  assign T_2289 = T_2286 | T_2288;
  assign GEN_59 = io_inner_release_bits_voluntary ? io_inner_release_bits_r_type : xact_vol_ir_r_type;
  assign GEN_60 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_id : xact_vol_ir_src;
  assign GEN_61 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_xact_id : xact_vol_ir_client_xact_id;
  assign T_2303 = T_2100 & T_2111;
  assign T_2307 = T_2303 ? 8'hff : 8'h0;
  assign T_2308 = ~ T_2307;
  assign T_2310 = 8'h1 << io_inner_release_bits_addr_beat;
  assign T_2311 = ~ T_2310;
  assign T_2312 = T_2308 | T_2311;
  assign T_2314 = T_2111 ? T_2312 : 8'h0;
  assign GEN_62 = T_2289 ? GEN_59 : xact_vol_ir_r_type;
  assign GEN_63 = T_2289 ? GEN_60 : xact_vol_ir_src;
  assign GEN_64 = T_2289 ? GEN_61 : xact_vol_ir_client_xact_id;
  assign GEN_65 = T_2289 ? T_2314 : GEN_57;
  assign T_2316 = T_2289 == 1'h0;
  assign T_2333 = pending_irel_data & T_2312;
  assign GEN_66 = T_2316 ? T_2333 : GEN_65;
  assign GEN_67 = T_2277 ? GEN_62 : xact_vol_ir_r_type;
  assign GEN_68 = T_2277 ? GEN_63 : xact_vol_ir_src;
  assign GEN_69 = T_2277 ? GEN_64 : xact_vol_ir_client_xact_id;
  assign GEN_70 = T_2277 ? GEN_66 : GEN_57;
  assign T_2334 = state == 4'h3;
  assign T_2335 = state == 4'h4;
  assign T_2337 = state == 4'h7;
  assign T_2338 = T_2334 | T_2335;
  assign T_2339 = T_2338 | T_2080;
  assign T_2340 = T_2339 | T_2337;
  assign T_2341 = T_2340 & vol_ignt_counter_pending;
  assign T_2343 = pending_irel_data != 8'h0;
  assign T_2344 = T_2343 | vol_ognt_counter_pending;
  assign T_2346 = T_2344 == 1'h0;
  assign T_2347 = T_2341 & T_2346;
  assign T_2379_addr_beat = 3'h0;
  assign T_2379_addr_block = xact_addr_block;
  assign T_2379_client_xact_id = xact_vol_ir_client_xact_id;
  assign T_2379_voluntary = 1'h1;
  assign T_2379_r_type = xact_vol_ir_r_type;
  assign T_2379_data = 64'h0;
  assign T_2379_client_id = xact_vol_ir_src;
  assign T_2440_addr_beat = 3'h0;
  assign T_2440_client_xact_id = T_2379_client_xact_id;
  assign T_2440_manager_xact_id = 2'h0;
  assign T_2440_is_builtin_type = 1'h1;
  assign T_2440_g_type = 4'h0;
  assign T_2440_data = 64'h0;
  assign T_2440_client_id = T_2379_client_id;
  assign GEN_0 = GEN_77;
  assign GEN_71 = 3'h1 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_72 = 3'h2 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_71;
  assign GEN_73 = 3'h3 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_72;
  assign GEN_74 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_73;
  assign GEN_75 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_74;
  assign GEN_76 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_75;
  assign GEN_77 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_76;
  assign T_2521 = GEN_0[0];
  assign GEN_1 = GEN_77;
  assign T_2522 = GEN_1[1];
  assign GEN_2 = GEN_77;
  assign T_2523 = GEN_2[2];
  assign GEN_3 = GEN_77;
  assign T_2524 = GEN_3[3];
  assign GEN_4 = GEN_77;
  assign T_2525 = GEN_4[4];
  assign GEN_5 = GEN_77;
  assign T_2526 = GEN_5[5];
  assign GEN_6 = GEN_77;
  assign T_2527 = GEN_6[6];
  assign GEN_7 = GEN_77;
  assign T_2528 = GEN_7[7];
  assign T_2532 = T_2521 ? 8'hff : 8'h0;
  assign T_2536 = T_2522 ? 8'hff : 8'h0;
  assign T_2540 = T_2523 ? 8'hff : 8'h0;
  assign T_2544 = T_2524 ? 8'hff : 8'h0;
  assign T_2548 = T_2525 ? 8'hff : 8'h0;
  assign T_2552 = T_2526 ? 8'hff : 8'h0;
  assign T_2556 = T_2527 ? 8'hff : 8'h0;
  assign T_2560 = T_2528 ? 8'hff : 8'h0;
  assign T_2561 = {T_2536,T_2532};
  assign T_2562 = {T_2544,T_2540};
  assign T_2563 = {T_2562,T_2561};
  assign T_2564 = {T_2552,T_2548};
  assign T_2565 = {T_2560,T_2556};
  assign T_2566 = {T_2565,T_2564};
  assign T_2567 = {T_2566,T_2563};
  assign T_2568 = ~ T_2567;
  assign T_2569 = T_2568 & io_inner_release_bits_data;
  assign GEN_8 = GEN_133;
  assign GEN_127 = 3'h1 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_128 = 3'h2 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_127;
  assign GEN_129 = 3'h3 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_128;
  assign GEN_130 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_129;
  assign GEN_131 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_130;
  assign GEN_132 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_131;
  assign GEN_133 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_132;
  assign T_2570 = T_2567 & GEN_8;
  assign T_2571 = T_2569 | T_2570;
  assign GEN_9 = T_2571;
  assign GEN_134 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_135 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_136 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_137 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_138 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_139 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_140 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_141 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_10 = 8'hff;
  assign GEN_142 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_0;
  assign GEN_143 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_1;
  assign GEN_144 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_2;
  assign GEN_145 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_3;
  assign GEN_146 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_4;
  assign GEN_147 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_5;
  assign GEN_148 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_6;
  assign GEN_149 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_7;
  assign GEN_160 = T_2303 ? GEN_134 : data_buffer_0;
  assign GEN_161 = T_2303 ? GEN_135 : data_buffer_1;
  assign GEN_162 = T_2303 ? GEN_136 : data_buffer_2;
  assign GEN_163 = T_2303 ? GEN_137 : data_buffer_3;
  assign GEN_164 = T_2303 ? GEN_138 : data_buffer_4;
  assign GEN_165 = T_2303 ? GEN_139 : data_buffer_5;
  assign GEN_166 = T_2303 ? GEN_140 : data_buffer_6;
  assign GEN_167 = T_2303 ? GEN_141 : data_buffer_7;
  assign GEN_169 = T_2303 ? GEN_142 : wmask_buffer_0;
  assign GEN_170 = T_2303 ? GEN_143 : wmask_buffer_1;
  assign GEN_171 = T_2303 ? GEN_144 : wmask_buffer_2;
  assign GEN_172 = T_2303 ? GEN_145 : wmask_buffer_3;
  assign GEN_173 = T_2303 ? GEN_146 : wmask_buffer_4;
  assign GEN_174 = T_2303 ? GEN_147 : wmask_buffer_5;
  assign GEN_175 = T_2303 ? GEN_148 : wmask_buffer_6;
  assign GEN_176 = T_2303 ? GEN_149 : wmask_buffer_7;
  assign T_2604_state = 2'h2;
  assign T_2631 = T_1653 | io_alloc_irel_should;
  assign T_2647 = T_2307 & T_2310;
  assign T_2648 = pending_orel_data | T_2647;
  assign T_2651 = io_outer_release_bits_r_type == 3'h0;
  assign T_2652 = io_outer_release_bits_r_type == 3'h1;
  assign T_2653 = io_outer_release_bits_r_type == 3'h2;
  assign T_2654 = T_2651 | T_2652;
  assign T_2655 = T_2654 | T_2653;
  assign T_2656 = T_2255 & T_2655;
  assign T_2660 = T_2656 ? 8'hff : 8'h0;
  assign T_2661 = ~ T_2660;
  assign T_2663 = 8'h1 << io_outer_release_bits_addr_beat;
  assign T_2664 = ~ T_2663;
  assign T_2665 = T_2661 | T_2664;
  assign T_2666 = T_2648 & T_2665;
  assign GEN_177 = T_2631 ? T_2666 : pending_orel_data;
  assign T_2677 = T_2655 == 1'h0;
  assign T_2679 = io_outer_release_bits_addr_beat == 3'h0;
  assign T_2680 = T_2677 | T_2679;
  assign GEN_179 = T_2680 ? 1'h1 : sending_orel;
  assign T_2692 = io_outer_release_bits_addr_beat == 3'h7;
  assign T_2693 = T_2677 | T_2692;
  assign GEN_180 = T_2693 ? 1'h0 : GEN_179;
  assign GEN_181 = T_2255 ? GEN_180 : sending_orel;
  assign GEN_182 = T_2255 ? 1'h0 : pending_orel_send;
  assign T_2702 = T_2255 & io_outer_release_bits_voluntary;
  assign T_2710 = T_2702 & T_2655;
  assign T_2714 = T_2712 == 3'h7;
  assign T_2716 = T_2712 + 3'h1;
  assign T_2717 = T_2716[2:0];
  assign GEN_183 = T_2710 ? T_2717 : T_2712;
  assign T_2718 = T_2710 & T_2714;
  assign T_2719 = T_2655 ? T_2712 : 3'h0;
  assign T_2720 = T_2655 ? T_2718 : T_2702;
  assign T_2723 = io_outer_grant_bits_g_type == 4'h0;
  assign T_2724 = io_outer_grant_bits_is_builtin_type & T_2723;
  assign T_2725 = T_2241 & T_2724;
  assign T_2733_0 = 3'h5;
  assign GEN_413 = {{1'd0}, T_2733_0};
  assign T_2735 = io_outer_grant_bits_g_type == GEN_413;
  assign T_2737 = io_outer_grant_bits_is_builtin_type ? T_2735 : T_2723;
  assign T_2739 = T_2725 & T_2737;
  assign T_2743 = T_2741 == 3'h7;
  assign T_2745 = T_2741 + 3'h1;
  assign T_2746 = T_2745[2:0];
  assign GEN_184 = T_2739 ? T_2746 : T_2741;
  assign T_2747 = T_2739 & T_2743;
  assign T_2748 = T_2737 ? T_2741 : 3'h0;
  assign T_2749 = T_2737 ? T_2747 : T_2725;
  assign T_2753 = T_2749 == 1'h0;
  assign T_2754 = T_2720 & T_2753;
  assign T_2756 = T_2751 + 1'h1;
  assign T_2757 = T_2756[0:0];
  assign GEN_185 = T_2754 ? T_2757 : T_2751;
  assign T_2759 = T_2720 == 1'h0;
  assign T_2760 = T_2749 & T_2759;
  assign T_2762 = T_2751 - 1'h1;
  assign T_2763 = T_2762[0:0];
  assign GEN_186 = T_2760 ? T_2763 : GEN_185;
  assign T_2765 = T_2751 > 1'h0;
  assign T_2774 = pending_orel_data >> vol_ognt_counter_up_idx;
  assign T_2775 = T_2774[0];
  assign T_2776 = T_2655 ? T_2775 : pending_orel_send;
  assign T_2777 = T_2337 & T_2776;
  assign T_2791 = T_2604_state == 2'h2;
  assign T_2792 = T_2791 ? 3'h0 : 3'h3;
  assign T_2828_addr_beat = vol_ognt_counter_up_idx;
  assign T_2828_addr_block = xact_addr_block;
  assign T_2828_client_xact_id = 2'h0;
  assign T_2828_voluntary = 1'h1;
  assign T_2828_r_type = T_2792;
  assign T_2828_data = GEN_11;
  assign GEN_11 = GEN_193;
  assign GEN_187 = 3'h1 == vol_ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_188 = 3'h2 == vol_ognt_counter_up_idx ? data_buffer_2 : GEN_187;
  assign GEN_189 = 3'h3 == vol_ognt_counter_up_idx ? data_buffer_3 : GEN_188;
  assign GEN_190 = 3'h4 == vol_ognt_counter_up_idx ? data_buffer_4 : GEN_189;
  assign GEN_191 = 3'h5 == vol_ognt_counter_up_idx ? data_buffer_5 : GEN_190;
  assign GEN_192 = 3'h6 == vol_ognt_counter_up_idx ? data_buffer_6 : GEN_191;
  assign GEN_193 = 3'h7 == vol_ognt_counter_up_idx ? data_buffer_7 : GEN_192;
  assign T_2857 = xact_iacq_is_builtin_type == 1'h0;
  assign T_2860 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_2871_0 = 3'h3;
  assign T_2873 = io_outer_acquire_bits_a_type == T_2871_0;
  assign T_2874 = io_outer_acquire_bits_is_builtin_type & T_2873;
  assign T_2875 = T_2860 & T_2874;
  assign T_2879 = T_2877 == 3'h7;
  assign T_2881 = T_2877 + 3'h1;
  assign T_2882 = T_2881[2:0];
  assign GEN_195 = T_2875 ? T_2882 : T_2877;
  assign T_2883 = T_2875 & T_2879;
  assign T_2884 = T_2874 ? T_2877 : xact_addr_beat;
  assign T_2885 = T_2874 ? T_2883 : T_2860;
  assign T_2891 = T_2724 == 1'h0;
  assign T_2892 = T_2241 & T_2891;
  assign T_2900_0 = 3'h5;
  assign GEN_414 = {{1'd0}, T_2900_0};
  assign T_2902 = io_outer_grant_bits_g_type == GEN_414;
  assign T_2904 = io_outer_grant_bits_is_builtin_type ? T_2902 : T_2723;
  assign T_2906 = T_2892 & T_2904;
  assign T_2910 = T_2908 == 3'h7;
  assign T_2912 = T_2908 + 3'h1;
  assign T_2913 = T_2912[2:0];
  assign GEN_196 = T_2906 ? T_2913 : T_2908;
  assign T_2914 = T_2906 & T_2910;
  assign T_2915 = T_2904 ? T_2908 : xact_addr_beat;
  assign T_2916 = T_2904 ? T_2914 : T_2892;
  assign T_2920 = T_2916 == 1'h0;
  assign T_2921 = T_2885 & T_2920;
  assign T_2923 = T_2918 + 1'h1;
  assign T_2924 = T_2923[0:0];
  assign GEN_197 = T_2921 ? T_2924 : T_2918;
  assign T_2926 = T_2885 == 1'h0;
  assign T_2927 = T_2916 & T_2926;
  assign T_2929 = T_2918 - 1'h1;
  assign T_2930 = T_2929[0:0];
  assign GEN_198 = T_2927 ? T_2930 : GEN_197;
  assign T_2932 = T_2918 > 1'h0;
  assign T_2933 = state == 4'h6;
  assign T_2937 = pending_put_data >> ognt_counter_up_idx;
  assign T_2938 = T_2937[0];
  assign T_2940 = T_2938 == 1'h0;
  assign T_2949_0 = 3'h2;
  assign T_2949_1 = 3'h3;
  assign T_2949_2 = 3'h4;
  assign T_2967 = xact_allocate | T_2940;
  assign T_2968 = T_2933 & T_2967;
  assign T_2971 = xact_op_code == 5'h1;
  assign T_2972 = xact_op_code == 5'h7;
  assign T_2973 = T_2971 | T_2972;
  assign T_2974 = xact_op_code[3];
  assign T_2975 = xact_op_code == 5'h4;
  assign T_2976 = T_2974 | T_2975;
  assign T_2977 = T_2973 | T_2976;
  assign T_2978 = xact_op_code == 5'h3;
  assign T_2979 = T_2977 | T_2978;
  assign T_2980 = xact_op_code == 5'h6;
  assign T_2981 = T_2979 | T_2980;
  assign T_2984 = {xact_op_code,1'h1};
  assign T_3015_addr_block = xact_addr_block;
  assign T_3015_client_xact_id = 2'h0;
  assign T_3015_addr_beat = 3'h0;
  assign T_3015_is_builtin_type = 1'h0;
  assign T_3015_a_type = {{2'd0}, T_2981};
  assign T_3015_union = {{5'd0}, T_2984};
  assign T_3015_data = 64'h0;
  assign GEN_12 = GEN_205;
  assign GEN_199 = 3'h1 == ognt_counter_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_200 = 3'h2 == ognt_counter_up_idx ? wmask_buffer_2 : GEN_199;
  assign GEN_201 = 3'h3 == ognt_counter_up_idx ? wmask_buffer_3 : GEN_200;
  assign GEN_202 = 3'h4 == ognt_counter_up_idx ? wmask_buffer_4 : GEN_201;
  assign GEN_203 = 3'h5 == ognt_counter_up_idx ? wmask_buffer_5 : GEN_202;
  assign GEN_204 = 3'h6 == ognt_counter_up_idx ? wmask_buffer_6 : GEN_203;
  assign GEN_205 = 3'h7 == ognt_counter_up_idx ? wmask_buffer_7 : GEN_204;
  assign T_3080 = {xact_op_code,1'h0};
  assign T_3081 = {xact_addr_byte,xact_op_size};
  assign T_3082 = {T_3081,T_3080};
  assign T_3084 = {xact_op_size,xact_op_code};
  assign T_3085 = {T_3084,1'h0};
  assign T_3087 = {GEN_12,1'h0};
  assign T_3099 = T_1993 ? 6'h2 : 6'h0;
  assign T_3101 = T_1995 ? 6'h0 : T_3099;
  assign T_3103 = T_1991 ? T_3082 : {{5'd0}, T_3101};
  assign T_3105 = T_2001 ? {{2'd0}, T_3087} : T_3103;
  assign T_3107 = T_1997 ? {{2'd0}, T_3087} : T_3105;
  assign T_3109 = T_2003 ? {{3'd0}, T_3085} : T_3107;
  assign T_3111 = T_1999 ? T_3082 : T_3109;
  assign T_3140_addr_block = xact_addr_block;
  assign T_3140_client_xact_id = 2'h0;
  assign T_3140_addr_beat = ognt_counter_up_idx;
  assign T_3140_is_builtin_type = 1'h1;
  assign T_3140_a_type = xact_iacq_a_type;
  assign T_3140_union = T_3111;
  assign T_3140_data = GEN_13;
  assign GEN_13 = GEN_212;
  assign GEN_206 = 3'h1 == ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_207 = 3'h2 == ognt_counter_up_idx ? data_buffer_2 : GEN_206;
  assign GEN_208 = 3'h3 == ognt_counter_up_idx ? data_buffer_3 : GEN_207;
  assign GEN_209 = 3'h4 == ognt_counter_up_idx ? data_buffer_4 : GEN_208;
  assign GEN_210 = 3'h5 == ognt_counter_up_idx ? data_buffer_5 : GEN_209;
  assign GEN_211 = 3'h6 == ognt_counter_up_idx ? data_buffer_6 : GEN_210;
  assign GEN_212 = 3'h7 == ognt_counter_up_idx ? data_buffer_7 : GEN_211;
  assign T_3168_addr_block = T_2857 ? T_3015_addr_block : T_3140_addr_block;
  assign T_3168_client_xact_id = T_2857 ? T_3015_client_xact_id : T_3140_client_xact_id;
  assign T_3168_addr_beat = T_2857 ? T_3015_addr_beat : T_3140_addr_beat;
  assign T_3168_is_builtin_type = T_2857 ? T_3015_is_builtin_type : T_3140_is_builtin_type;
  assign T_3168_a_type = T_2857 ? T_3015_a_type : T_3140_a_type;
  assign T_3168_union = T_2857 ? T_3015_union : T_3140_union;
  assign T_3168_data = T_2857 ? T_3015_data : T_3140_data;
  assign T_3197 = T_2933 & ognt_counter_up_done;
  assign GEN_213 = T_3197 ? 4'h7 : GEN_58;
  assign GEN_214 = ognt_counter_pending ? 1'h1 : vol_ognt_counter_pending;
  assign T_3207_0 = 3'h5;
  assign T_3207_1 = 3'h4;
  assign GEN_415 = {{1'd0}, T_3207_0};
  assign T_3209 = io_outer_grant_bits_g_type == GEN_415;
  assign GEN_416 = {{1'd0}, T_3207_1};
  assign T_3210 = io_outer_grant_bits_g_type == GEN_416;
  assign T_3211 = T_3209 | T_3210;
  assign T_3213 = io_outer_grant_bits_is_builtin_type ? T_3211 : T_2723;
  assign T_3214 = T_2241 & T_3213;
  assign GEN_14 = GEN_221;
  assign GEN_215 = 3'h1 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_216 = 3'h2 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_215;
  assign GEN_217 = 3'h3 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_216;
  assign GEN_218 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_217;
  assign GEN_219 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_218;
  assign GEN_220 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_219;
  assign GEN_221 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_220;
  assign T_3215 = GEN_14[0];
  assign GEN_15 = GEN_221;
  assign T_3216 = GEN_15[1];
  assign GEN_16 = GEN_221;
  assign T_3217 = GEN_16[2];
  assign GEN_17 = GEN_221;
  assign T_3218 = GEN_17[3];
  assign GEN_18 = GEN_221;
  assign T_3219 = GEN_18[4];
  assign GEN_19 = GEN_221;
  assign T_3220 = GEN_19[5];
  assign GEN_20 = GEN_221;
  assign T_3221 = GEN_20[6];
  assign GEN_21 = GEN_221;
  assign T_3222 = GEN_21[7];
  assign T_3226 = T_3215 ? 8'hff : 8'h0;
  assign T_3230 = T_3216 ? 8'hff : 8'h0;
  assign T_3234 = T_3217 ? 8'hff : 8'h0;
  assign T_3238 = T_3218 ? 8'hff : 8'h0;
  assign T_3242 = T_3219 ? 8'hff : 8'h0;
  assign T_3246 = T_3220 ? 8'hff : 8'h0;
  assign T_3250 = T_3221 ? 8'hff : 8'h0;
  assign T_3254 = T_3222 ? 8'hff : 8'h0;
  assign T_3255 = {T_3230,T_3226};
  assign T_3256 = {T_3238,T_3234};
  assign T_3257 = {T_3256,T_3255};
  assign T_3258 = {T_3246,T_3242};
  assign T_3259 = {T_3254,T_3250};
  assign T_3260 = {T_3259,T_3258};
  assign T_3261 = {T_3260,T_3257};
  assign T_3262 = ~ T_3261;
  assign T_3263 = T_3262 & io_outer_grant_bits_data;
  assign GEN_22 = GEN_277;
  assign GEN_271 = 3'h1 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_272 = 3'h2 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_271;
  assign GEN_273 = 3'h3 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_272;
  assign GEN_274 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_273;
  assign GEN_275 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_274;
  assign GEN_276 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_275;
  assign GEN_277 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_276;
  assign T_3264 = T_3261 & GEN_22;
  assign T_3265 = T_3263 | T_3264;
  assign GEN_23 = T_3265;
  assign GEN_278 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_160;
  assign GEN_279 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_161;
  assign GEN_280 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_162;
  assign GEN_281 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_163;
  assign GEN_282 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_164;
  assign GEN_283 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_165;
  assign GEN_284 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_166;
  assign GEN_285 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_167;
  assign GEN_24 = 8'hff;
  assign GEN_286 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_169;
  assign GEN_287 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_170;
  assign GEN_288 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_171;
  assign GEN_289 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_172;
  assign GEN_290 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_173;
  assign GEN_291 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_174;
  assign GEN_292 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_175;
  assign GEN_293 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_176;
  assign GEN_304 = T_3214 ? GEN_278 : GEN_160;
  assign GEN_305 = T_3214 ? GEN_279 : GEN_161;
  assign GEN_306 = T_3214 ? GEN_280 : GEN_162;
  assign GEN_307 = T_3214 ? GEN_281 : GEN_163;
  assign GEN_308 = T_3214 ? GEN_282 : GEN_164;
  assign GEN_309 = T_3214 ? GEN_283 : GEN_165;
  assign GEN_310 = T_3214 ? GEN_284 : GEN_166;
  assign GEN_311 = T_3214 ? GEN_285 : GEN_167;
  assign GEN_313 = T_3214 ? GEN_286 : GEN_169;
  assign GEN_314 = T_3214 ? GEN_287 : GEN_170;
  assign GEN_315 = T_3214 ? GEN_288 : GEN_171;
  assign GEN_316 = T_3214 ? GEN_289 : GEN_172;
  assign GEN_317 = T_3214 ? GEN_290 : GEN_173;
  assign GEN_318 = T_3214 ? GEN_291 : GEN_174;
  assign GEN_319 = T_3214 ? GEN_292 : GEN_175;
  assign GEN_320 = T_3214 ? GEN_293 : GEN_176;
  assign T_3268 = scoreboard_3 | ognt_counter_pending;
  assign T_3269 = T_3268 | vol_ognt_counter_pending;
  assign T_3281 = T_2179 == 1'h0;
  assign T_3283 = T_2175 & T_3281;
  assign T_3291_0 = 3'h5;
  assign GEN_417 = {{1'd0}, T_3291_0};
  assign T_3293 = io_inner_grant_bits_g_type == GEN_417;
  assign T_3295 = io_inner_grant_bits_is_builtin_type ? T_3293 : T_2178;
  assign T_3297 = T_3283 & T_3295;
  assign T_3301 = T_3299 == 3'h7;
  assign T_3303 = T_3299 + 3'h1;
  assign T_3304 = T_3303[2:0];
  assign GEN_321 = T_3297 ? T_3304 : T_3299;
  assign T_3305 = T_3297 & T_3301;
  assign T_3306 = T_3295 ? T_3299 : 3'h0;
  assign T_3307 = T_3295 ? T_3305 : T_3283;
  assign T_3308 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3326 = T_3308 == 1'h0;
  assign T_3327 = T_3307 & T_3326;
  assign T_3329 = T_3324 + 1'h1;
  assign T_3330 = T_3329[0:0];
  assign GEN_323 = T_3327 ? T_3330 : T_3324;
  assign T_3332 = T_3307 == 1'h0;
  assign T_3333 = T_3308 & T_3332;
  assign T_3335 = T_3324 - 1'h1;
  assign T_3336 = T_3335[0:0];
  assign GEN_324 = T_3333 ? T_3336 : GEN_323;
  assign T_3338 = T_3324 > 1'h0;
  assign T_3343 = T_1798 == 1'h0;
  assign T_3360 = pending_ignt_data | T_2647;
  assign T_3370_0 = 3'h5;
  assign T_3370_1 = 3'h4;
  assign GEN_418 = {{1'd0}, T_3370_0};
  assign T_3372 = io_outer_grant_bits_g_type == GEN_418;
  assign GEN_419 = {{1'd0}, T_3370_1};
  assign T_3373 = io_outer_grant_bits_g_type == GEN_419;
  assign T_3374 = T_3372 | T_3373;
  assign T_3376 = io_outer_grant_bits_is_builtin_type ? T_3374 : T_2723;
  assign T_3377 = T_2241 & T_3376;
  assign T_3382 = T_3377 ? 8'hff : 8'h0;
  assign T_3384 = 8'h1 << io_outer_grant_bits_addr_beat;
  assign T_3385 = T_3382 & T_3384;
  assign T_3386 = T_3360 | T_3385;
  assign GEN_327 = T_3343 ? T_3386 : GEN_45;
  assign T_3389 = state == 4'h1;
  assign T_3390 = T_1611 | T_3389;
  assign T_3393 = T_3390 | scoreboard_0;
  assign T_3395 = T_3393 == 1'h0;
  assign T_3412 = 3'h6 == ignt_q_io_deq_bits_a_type;
  assign T_3413 = T_3412 ? 3'h1 : 3'h3;
  assign T_3414 = 3'h5 == ignt_q_io_deq_bits_a_type;
  assign T_3415 = T_3414 ? 3'h1 : T_3413;
  assign T_3416 = 3'h4 == ignt_q_io_deq_bits_a_type;
  assign T_3417 = T_3416 ? 3'h4 : T_3415;
  assign T_3418 = 3'h3 == ignt_q_io_deq_bits_a_type;
  assign T_3419 = T_3418 ? 3'h3 : T_3417;
  assign T_3420 = 3'h2 == ignt_q_io_deq_bits_a_type;
  assign T_3421 = T_3420 ? 3'h3 : T_3419;
  assign T_3422 = 3'h1 == ignt_q_io_deq_bits_a_type;
  assign T_3423 = T_3422 ? 3'h5 : T_3421;
  assign T_3424 = 3'h0 == ignt_q_io_deq_bits_a_type;
  assign T_3425 = T_3424 ? 3'h4 : T_3423;
  assign T_3426 = ignt_q_io_deq_bits_is_builtin_type ? T_3425 : 3'h0;
  assign T_3455_addr_beat = ignt_q_io_deq_bits_addr_beat;
  assign T_3455_client_xact_id = ignt_q_io_deq_bits_client_xact_id;
  assign T_3455_manager_xact_id = 2'h2;
  assign T_3455_is_builtin_type = ignt_q_io_deq_bits_is_builtin_type;
  assign T_3455_g_type = {{1'd0}, T_3426};
  assign T_3455_data = GEN_25;
  assign T_3455_client_id = ignt_q_io_deq_bits_client_id;
  assign GEN_25 = GEN_334;
  assign GEN_328 = 3'h1 == ignt_data_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_329 = 3'h2 == ignt_data_idx ? data_buffer_2 : GEN_328;
  assign GEN_330 = 3'h3 == ignt_data_idx ? data_buffer_3 : GEN_329;
  assign GEN_331 = 3'h4 == ignt_data_idx ? data_buffer_4 : GEN_330;
  assign GEN_332 = 3'h5 == ignt_data_idx ? data_buffer_5 : GEN_331;
  assign GEN_333 = 3'h6 == ignt_data_idx ? data_buffer_6 : GEN_332;
  assign GEN_334 = 3'h7 == ignt_data_idx ? data_buffer_7 : GEN_333;
  assign T_3491_0 = 3'h5;
  assign GEN_420 = {{1'd0}, T_3491_0};
  assign T_3493 = io_inner_grant_bits_g_type == GEN_420;
  assign T_3495 = io_inner_grant_bits_is_builtin_type ? T_3493 : T_2178;
  assign T_3497 = T_2175 & T_3495;
  assign T_3501 = T_3499 == 3'h7;
  assign T_3503 = T_3499 + 3'h1;
  assign T_3504 = T_3503[2:0];
  assign GEN_335 = T_3497 ? T_3504 : T_3499;
  assign T_3505 = T_3497 & T_3501;
  assign T_3506 = T_3495 ? T_3499 : ignt_q_io_deq_bits_addr_beat;
  assign T_3507 = T_3495 ? T_3505 : T_2175;
  assign T_3512 = T_2337 & scoreboard_6;
  assign T_3514 = T_3269 == 1'h0;
  assign T_3522_0 = 3'h5;
  assign T_3522_1 = 3'h4;
  assign GEN_421 = {{1'd0}, T_3522_0};
  assign T_3524 = io_inner_grant_bits_g_type == GEN_421;
  assign GEN_422 = {{1'd0}, T_3522_1};
  assign T_3525 = io_inner_grant_bits_g_type == GEN_422;
  assign T_3526 = T_3524 | T_3525;
  assign T_3528 = io_inner_grant_bits_is_builtin_type ? T_3526 : T_2178;
  assign T_3529 = pending_ignt_data >> ignt_data_idx;
  assign T_3530 = T_3529[0];
  assign T_3532 = T_3528 ? T_3530 : T_3395;
  assign T_3533 = T_3514 & T_3532;
  assign GEN_338 = T_3512 ? T_3533 : T_2347;
  assign GEN_339 = T_2250 ? ignt_data_done : 1'h0;
  assign GEN_340 = T_2250 ? ignt_data_idx : T_2440_addr_beat;
  assign GEN_341 = T_2250 ? T_3455_client_xact_id : T_2440_client_xact_id;
  assign GEN_342 = T_2250 ? T_3455_manager_xact_id : T_2440_manager_xact_id;
  assign GEN_343 = T_2250 ? T_3455_is_builtin_type : T_2440_is_builtin_type;
  assign GEN_344 = T_2250 ? T_3455_g_type : T_2440_g_type;
  assign GEN_345 = T_2250 ? T_3455_data : T_2440_data;
  assign GEN_346 = T_2250 ? T_3455_client_id : T_2440_client_id;
  assign GEN_349 = T_2250 ? GEN_338 : T_2347;
  assign T_3540 = ~ io_incoherent_0;
  assign GEN_350 = T_1798 ? {{1'd0}, T_3540} : T_2079;
  assign T_3551 = T_1767 & io_inner_acquire_valid;
  assign T_3552 = T_1798 | T_3551;
  assign T_3562_0 = 3'h2;
  assign T_3562_1 = 3'h3;
  assign T_3562_2 = 3'h4;
  assign T_3564 = io_inner_acquire_bits_a_type == T_3562_0;
  assign T_3565 = io_inner_acquire_bits_a_type == T_3562_1;
  assign T_3566 = io_inner_acquire_bits_a_type == T_3562_2;
  assign T_3567 = T_3564 | T_3565;
  assign T_3568 = T_3567 | T_3566;
  assign T_3569 = io_inner_acquire_bits_is_builtin_type & T_3568;
  assign T_3570 = T_1612 & T_3569;
  assign T_3571 = T_3570 & T_3552;
  assign T_3573 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3574 = io_inner_acquire_bits_is_builtin_type & T_3573;
  assign T_3603 = T_1921 | T_1918;
  assign T_3604 = io_inner_acquire_bits_union[8:1];
  assign T_3606 = T_3603 ? T_3604 : 8'h0;
  assign T_3607 = T_3574 ? 8'hff : T_3606;
  assign T_3608 = T_3607[0];
  assign T_3609 = T_3607[1];
  assign T_3610 = T_3607[2];
  assign T_3611 = T_3607[3];
  assign T_3612 = T_3607[4];
  assign T_3613 = T_3607[5];
  assign T_3614 = T_3607[6];
  assign T_3615 = T_3607[7];
  assign T_3619 = T_3608 ? 8'hff : 8'h0;
  assign T_3623 = T_3609 ? 8'hff : 8'h0;
  assign T_3627 = T_3610 ? 8'hff : 8'h0;
  assign T_3631 = T_3611 ? 8'hff : 8'h0;
  assign T_3635 = T_3612 ? 8'hff : 8'h0;
  assign T_3639 = T_3613 ? 8'hff : 8'h0;
  assign T_3643 = T_3614 ? 8'hff : 8'h0;
  assign T_3647 = T_3615 ? 8'hff : 8'h0;
  assign T_3648 = {T_3623,T_3619};
  assign T_3649 = {T_3631,T_3627};
  assign T_3650 = {T_3649,T_3648};
  assign T_3651 = {T_3639,T_3635};
  assign T_3652 = {T_3647,T_3643};
  assign T_3653 = {T_3652,T_3651};
  assign T_3654 = {T_3653,T_3650};
  assign T_3655 = ~ T_3654;
  assign GEN_26 = GEN_357;
  assign GEN_351 = 3'h1 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_352 = 3'h2 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_351;
  assign GEN_353 = 3'h3 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_352;
  assign GEN_354 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_353;
  assign GEN_355 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_354;
  assign GEN_356 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_355;
  assign GEN_357 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_356;
  assign T_3656 = T_3655 & GEN_26;
  assign T_3657 = T_3654 & io_inner_acquire_bits_data;
  assign T_3658 = T_3656 | T_3657;
  assign GEN_27 = T_3658;
  assign GEN_358 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_304;
  assign GEN_359 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_305;
  assign GEN_360 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_306;
  assign GEN_361 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_307;
  assign GEN_362 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_308;
  assign GEN_363 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_309;
  assign GEN_364 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_310;
  assign GEN_365 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_311;
  assign GEN_28 = GEN_372;
  assign GEN_366 = 3'h1 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_367 = 3'h2 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_366;
  assign GEN_368 = 3'h3 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_367;
  assign GEN_369 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_368;
  assign GEN_370 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_369;
  assign GEN_371 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_370;
  assign GEN_372 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_371;
  assign T_3695 = T_3607 | GEN_28;
  assign GEN_29 = T_3695;
  assign GEN_373 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_313;
  assign GEN_374 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_314;
  assign GEN_375 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_315;
  assign GEN_376 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_316;
  assign GEN_377 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_317;
  assign GEN_378 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_318;
  assign GEN_379 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_319;
  assign GEN_380 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_320;
  assign GEN_383 = T_3571 ? GEN_358 : GEN_304;
  assign GEN_384 = T_3571 ? GEN_359 : GEN_305;
  assign GEN_385 = T_3571 ? GEN_360 : GEN_306;
  assign GEN_386 = T_3571 ? GEN_361 : GEN_307;
  assign GEN_387 = T_3571 ? GEN_362 : GEN_308;
  assign GEN_388 = T_3571 ? GEN_363 : GEN_309;
  assign GEN_389 = T_3571 ? GEN_364 : GEN_310;
  assign GEN_390 = T_3571 ? GEN_365 : GEN_311;
  assign GEN_393 = T_3571 ? GEN_373 : GEN_313;
  assign GEN_394 = T_3571 ? GEN_374 : GEN_314;
  assign GEN_395 = T_3571 ? GEN_375 : GEN_315;
  assign GEN_396 = T_3571 ? GEN_376 : GEN_316;
  assign GEN_397 = T_3571 ? GEN_377 : GEN_317;
  assign GEN_398 = T_3571 ? GEN_378 : GEN_318;
  assign GEN_399 = T_3571 ? GEN_379 : GEN_319;
  assign GEN_400 = T_3571 ? GEN_380 : GEN_320;
  assign T_3698 = scoreboard_0 | T_2343;
  assign T_3699 = T_3698 | vol_ignt_counter_pending;
  assign T_3700 = T_3699 | scoreboard_3;
  assign T_3701 = T_3700 | vol_ognt_counter_pending;
  assign T_3702 = T_3701 | ognt_counter_pending;
  assign T_3703 = T_3702 | scoreboard_6;
  assign T_3704 = T_3703 | ifin_counter_pending;
  assign T_3706 = T_3704 == 1'h0;
  assign T_3708 = T_2337 & all_pending_done;
  assign GEN_401 = T_3708 ? 4'h0 : GEN_213;
  assign GEN_402 = T_3708 ? 8'h0 : GEN_393;
  assign GEN_403 = T_3708 ? 8'h0 : GEN_394;
  assign GEN_404 = T_3708 ? 8'h0 : GEN_395;
  assign GEN_405 = T_3708 ? 8'h0 : GEN_396;
  assign GEN_406 = T_3708 ? 8'h0 : GEN_397;
  assign GEN_407 = T_3708 ? 8'h0 : GEN_398;
  assign GEN_408 = T_3708 ? 8'h0 : GEN_399;
  assign GEN_409 = T_3708 ? 8'h0 : GEN_400;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_121[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_122[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  state = GEN_32[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  xact_addr_block = GEN_33[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  xact_allocate = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  xact_amo_shift_bytes = GEN_42[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  xact_op_code = GEN_43[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  xact_addr_byte = GEN_47[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_78 = {1{$random}};
  xact_op_size = GEN_78[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_79 = {1{$random}};
  xact_vol_ir_r_type = GEN_79[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_80 = {1{$random}};
  xact_vol_ir_src = GEN_80[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_81 = {1{$random}};
  xact_vol_ir_client_xact_id = GEN_81[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_82 = {1{$random}};
  pending_irel_data = GEN_82[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_83 = {1{$random}};
  pending_put_data = GEN_83[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_84 = {1{$random}};
  pending_ignt_data = GEN_84[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {1{$random}};
  pending_iprbs = GEN_85[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  pending_orel_send = GEN_86[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_87 = {1{$random}};
  pending_orel_data = GEN_87[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  sending_orel = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {2{$random}};
  data_buffer_0 = GEN_89[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {2{$random}};
  data_buffer_1 = GEN_90[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {2{$random}};
  data_buffer_2 = GEN_91[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_92 = {2{$random}};
  data_buffer_3 = GEN_92[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_93 = {2{$random}};
  data_buffer_4 = GEN_93[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_94 = {2{$random}};
  data_buffer_5 = GEN_94[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_95 = {2{$random}};
  data_buffer_6 = GEN_95[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_96 = {2{$random}};
  data_buffer_7 = GEN_96[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_97 = {1{$random}};
  wmask_buffer_0 = GEN_97[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_98 = {1{$random}};
  wmask_buffer_1 = GEN_98[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_99 = {1{$random}};
  wmask_buffer_2 = GEN_99[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {1{$random}};
  wmask_buffer_3 = GEN_100[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_101 = {1{$random}};
  wmask_buffer_4 = GEN_101[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_102 = {1{$random}};
  wmask_buffer_5 = GEN_102[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_103 = {1{$random}};
  wmask_buffer_6 = GEN_103[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_104 = {1{$random}};
  wmask_buffer_7 = GEN_104[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_105 = {1{$random}};
  T_2091 = GEN_105[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_106 = {1{$random}};
  T_2115 = GEN_106[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_107 = {1{$random}};
  T_2125 = GEN_107[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_108 = {1{$random}};
  T_2166 = GEN_108[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_109 = {1{$random}};
  T_2197 = GEN_109[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_110 = {1{$random}};
  T_2207 = GEN_110[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_111 = {1{$random}};
  T_2712 = GEN_111[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {1{$random}};
  T_2741 = GEN_112[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_113 = {1{$random}};
  T_2751 = GEN_113[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_114 = {1{$random}};
  T_2877 = GEN_114[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  T_2908 = GEN_115[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_116 = {1{$random}};
  T_2918 = GEN_116[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_117 = {1{$random}};
  T_3299 = GEN_117[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_118 = {1{$random}};
  T_3314 = GEN_118[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  T_3324 = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  T_3499 = GEN_120[2:0];
  `endif
  GEN_121 = {1{$random}};
  GEN_122 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_3708) begin
        state <= 4'h0;
      end else begin
        if(T_3197) begin
          state <= 4'h7;
        end else begin
          if(T_2224) begin
            state <= 4'h7;
          end else begin
            if(T_2146) begin
              if(T_2055) begin
                state <= 4'h6;
              end else begin
                state <= 4'h7;
              end
            end else begin
              if(T_1798) begin
                state <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      xact_addr_block <= 26'h0;
    end else begin
      if(T_2224) begin
        xact_addr_block <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1798) begin
          xact_addr_block <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_allocate <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_amo_shift_bytes <= T_1915;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        if(T_1922) begin
          xact_op_code <= 5'h1;
        end else begin
          xact_op_code <= T_1923;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_addr_byte <= T_1925;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_op_size <= T_1926;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_r_type <= io_inner_release_bits_r_type;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_src <= io_inner_release_bits_client_id;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_client_xact_id <= io_inner_release_bits_client_xact_id;
          end
        end
      end
    end
    if(reset) begin
      pending_irel_data <= 8'h0;
    end else begin
      if(T_2277) begin
        if(T_2316) begin
          pending_irel_data <= T_2333;
        end else begin
          if(T_2289) begin
            if(T_2111) begin
              pending_irel_data <= T_2312;
            end else begin
              pending_irel_data <= 8'h0;
            end
          end else begin
            if(T_2224) begin
              pending_irel_data <= 8'hff;
            end
          end
        end
      end else begin
        if(T_2224) begin
          pending_irel_data <= 8'hff;
        end
      end
    end
    if(reset) begin
      pending_put_data <= 8'h0;
    end else begin
      if(T_1798) begin
        if(T_1921) begin
          pending_put_data <= T_1956;
        end else begin
          pending_put_data <= 8'h0;
        end
      end else begin
        if(T_1852) begin
          pending_put_data <= T_1907;
        end
      end
    end
    if(reset) begin
      pending_ignt_data <= 8'h0;
    end else begin
      if(T_3343) begin
        pending_ignt_data <= T_3386;
      end else begin
        if(T_1798) begin
          pending_ignt_data <= 8'h0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      pending_iprbs <= GEN_350[0];
    end
    if(reset) begin
      pending_orel_send <= 1'h0;
    end else begin
      if(T_2255) begin
        pending_orel_send <= 1'h0;
      end
    end
    if(reset) begin
      pending_orel_data <= 8'h0;
    end else begin
      if(T_2631) begin
        pending_orel_data <= T_2666;
      end
    end
    if(reset) begin
      sending_orel <= 1'h0;
    end else begin
      if(T_2255) begin
        if(T_2693) begin
          sending_orel <= 1'h0;
        end else begin
          if(T_2680) begin
            sending_orel <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1691_0;
    end else begin
      if(T_3571) begin
        if(3'h0 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h0 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h0 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1691_1;
    end else begin
      if(T_3571) begin
        if(3'h1 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h1 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h1 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1691_2;
    end else begin
      if(T_3571) begin
        if(3'h2 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h2 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h2 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1691_3;
    end else begin
      if(T_3571) begin
        if(3'h3 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h3 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h3 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1691_4;
    end else begin
      if(T_3571) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1691_5;
    end else begin
      if(T_3571) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1691_6;
    end else begin
      if(T_3571) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1691_7;
    end else begin
      if(T_3571) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1709_0;
    end else begin
      if(T_3708) begin
        wmask_buffer_0 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h0 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h0 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h0 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_0 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_0 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1709_1;
    end else begin
      if(T_3708) begin
        wmask_buffer_1 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h1 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h1 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h1 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_1 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_1 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1709_2;
    end else begin
      if(T_3708) begin
        wmask_buffer_2 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h2 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h2 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h2 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_2 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_2 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1709_3;
    end else begin
      if(T_3708) begin
        wmask_buffer_3 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h3 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h3 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h3 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_3 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_3 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1709_4;
    end else begin
      if(T_3708) begin
        wmask_buffer_4 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h4 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h4 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_4 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_4 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1709_5;
    end else begin
      if(T_3708) begin
        wmask_buffer_5 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h5 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h5 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_5 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_5 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1709_6;
    end else begin
      if(T_3708) begin
        wmask_buffer_6 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h6 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h6 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_6 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_6 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1709_7;
    end else begin
      if(T_3708) begin
        wmask_buffer_7 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h7 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h7 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_7 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_7 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_2091 <= 3'h0;
    end
    if(reset) begin
      T_2115 <= 3'h0;
    end else begin
      if(T_2113) begin
        T_2115 <= T_2120;
      end
    end
    if(reset) begin
      T_2125 <= 1'h0;
    end else begin
      if(T_2134) begin
        T_2125 <= T_2137;
      end else begin
        if(T_2128) begin
          T_2125 <= T_2131;
        end
      end
    end
    if(reset) begin
      T_2166 <= 3'h0;
    end else begin
      if(T_2164) begin
        T_2166 <= T_2171;
      end
    end
    if(reset) begin
      T_2197 <= 3'h0;
    end else begin
      if(T_2195) begin
        T_2197 <= T_2202;
      end
    end
    if(reset) begin
      T_2207 <= 1'h0;
    end else begin
      if(T_2216) begin
        T_2207 <= T_2219;
      end else begin
        if(T_2210) begin
          T_2207 <= T_2213;
        end
      end
    end
    if(reset) begin
      T_2712 <= 3'h0;
    end else begin
      if(T_2710) begin
        T_2712 <= T_2717;
      end
    end
    if(reset) begin
      T_2741 <= 3'h0;
    end else begin
      if(T_2739) begin
        T_2741 <= T_2746;
      end
    end
    if(reset) begin
      T_2751 <= 1'h0;
    end else begin
      if(T_2760) begin
        T_2751 <= T_2763;
      end else begin
        if(T_2754) begin
          T_2751 <= T_2757;
        end
      end
    end
    if(reset) begin
      T_2877 <= 3'h0;
    end else begin
      if(T_2875) begin
        T_2877 <= T_2882;
      end
    end
    if(reset) begin
      T_2908 <= 3'h0;
    end else begin
      if(T_2906) begin
        T_2908 <= T_2913;
      end
    end
    if(reset) begin
      T_2918 <= 1'h0;
    end else begin
      if(T_2927) begin
        T_2918 <= T_2930;
      end else begin
        if(T_2921) begin
          T_2918 <= T_2924;
        end
      end
    end
    if(reset) begin
      T_3299 <= 3'h0;
    end else begin
      if(T_3297) begin
        T_3299 <= T_3304;
      end
    end
    if(reset) begin
      T_3314 <= 3'h0;
    end
    if(reset) begin
      T_3324 <= 1'h0;
    end else begin
      if(T_3333) begin
        T_3324 <= T_3336;
      end else begin
        if(T_3327) begin
          T_3324 <= T_3330;
        end
      end
    end
    if(reset) begin
      T_3499 <= 3'h0;
    end else begin
      if(T_3497) begin
        T_3499 <= T_3504;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1652) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:98 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1652) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1666) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1677) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:105 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1677) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module LockingRRArbiter_5(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [10:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [10:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [1:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_addr_beat,
  input   io_in_2_bits_is_builtin_type,
  input  [2:0] io_in_2_bits_a_type,
  input  [10:0] io_in_2_bits_union,
  input  [63:0] io_in_2_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [10:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [25:0] GEN_0_bits_addr_block;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire [2:0] GEN_0_bits_addr_beat;
  wire  GEN_0_bits_is_builtin_type;
  wire [2:0] GEN_0_bits_a_type;
  wire [10:0] GEN_0_bits_union;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_8;
  wire  GEN_9;
  wire [25:0] GEN_10;
  wire [1:0] GEN_11;
  wire [2:0] GEN_12;
  wire  GEN_13;
  wire [2:0] GEN_14;
  wire [10:0] GEN_15;
  wire [63:0] GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [25:0] GEN_19;
  wire [1:0] GEN_20;
  wire [2:0] GEN_21;
  wire  GEN_22;
  wire [2:0] GEN_23;
  wire [10:0] GEN_24;
  wire [63:0] GEN_25;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [25:0] GEN_1_bits_addr_block;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire [2:0] GEN_1_bits_addr_beat;
  wire  GEN_1_bits_is_builtin_type;
  wire [2:0] GEN_1_bits_a_type;
  wire [10:0] GEN_1_bits_union;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [25:0] GEN_2_bits_addr_block;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire [2:0] GEN_2_bits_addr_beat;
  wire  GEN_2_bits_is_builtin_type;
  wire [2:0] GEN_2_bits_a_type;
  wire [10:0] GEN_2_bits_union;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [25:0] GEN_3_bits_addr_block;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire [2:0] GEN_3_bits_addr_beat;
  wire  GEN_3_bits_is_builtin_type;
  wire [2:0] GEN_3_bits_a_type;
  wire [10:0] GEN_3_bits_union;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [25:0] GEN_4_bits_addr_block;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire [2:0] GEN_4_bits_addr_beat;
  wire  GEN_4_bits_is_builtin_type;
  wire [2:0] GEN_4_bits_a_type;
  wire [10:0] GEN_4_bits_union;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [25:0] GEN_5_bits_addr_block;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire [2:0] GEN_5_bits_addr_beat;
  wire  GEN_5_bits_is_builtin_type;
  wire [2:0] GEN_5_bits_a_type;
  wire [10:0] GEN_5_bits_union;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [25:0] GEN_6_bits_addr_block;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire [2:0] GEN_6_bits_addr_beat;
  wire  GEN_6_bits_is_builtin_type;
  wire [2:0] GEN_6_bits_a_type;
  wire [10:0] GEN_6_bits_union;
  wire [63:0] GEN_6_bits_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [25:0] GEN_7_bits_addr_block;
  wire [1:0] GEN_7_bits_client_xact_id;
  wire [2:0] GEN_7_bits_addr_beat;
  wire  GEN_7_bits_is_builtin_type;
  wire [2:0] GEN_7_bits_a_type;
  wire [10:0] GEN_7_bits_union;
  wire [63:0] GEN_7_bits_data;
  reg [2:0] T_882;
  reg [31:0] GEN_0;
  reg [1:0] T_884;
  reg [31:0] GEN_1;
  wire  T_886;
  wire [2:0] T_895_0;
  wire  T_897;
  wire  T_898;
  wire  T_899;
  wire  T_900;
  wire [3:0] T_904;
  wire [2:0] T_905;
  wire [1:0] GEN_152;
  wire [2:0] GEN_153;
  wire [1:0] GEN_154;
  reg [1:0] lastGrant;
  reg [31:0] GEN_2;
  wire [1:0] GEN_155;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  validMask_1;
  wire  validMask_2;
  wire  T_912;
  wire  T_913;
  wire  T_914;
  wire  T_918;
  wire  T_920;
  wire  T_922;
  wire  T_924;
  wire  T_928;
  wire  T_929;
  wire  T_930;
  wire  T_932;
  wire  T_933;
  wire  T_934;
  wire  T_936;
  wire  T_937;
  wire  T_938;
  wire  T_940;
  wire  T_941;
  wire  T_942;
  wire [1:0] GEN_156;
  wire [1:0] GEN_157;
  wire [1:0] GEN_158;
  wire [1:0] GEN_159;
  assign io_in_0_ready = T_934;
  assign io_in_1_ready = T_938;
  assign io_in_2_ready = T_942;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_block = GEN_1_bits_addr_block;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_addr_beat = GEN_3_bits_addr_beat;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_a_type = GEN_5_bits_a_type;
  assign io_out_bits_union = GEN_6_bits_union;
  assign io_out_bits_data = GEN_7_bits_data;
  assign io_chosen = GEN_154;
  assign choice = GEN_159;
  assign GEN_0_ready = GEN_17;
  assign GEN_0_valid = GEN_18;
  assign GEN_0_bits_addr_block = GEN_19;
  assign GEN_0_bits_client_xact_id = GEN_20;
  assign GEN_0_bits_addr_beat = GEN_21;
  assign GEN_0_bits_is_builtin_type = GEN_22;
  assign GEN_0_bits_a_type = GEN_23;
  assign GEN_0_bits_union = GEN_24;
  assign GEN_0_bits_data = GEN_25;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_ready : GEN_8;
  assign GEN_18 = 2'h2 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_addr_block : GEN_10;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_11;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_12;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_13;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_a_type : GEN_14;
  assign GEN_24 = 2'h2 == io_chosen ? io_in_2_bits_union : GEN_15;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_data : GEN_16;
  assign GEN_1_ready = GEN_17;
  assign GEN_1_valid = GEN_18;
  assign GEN_1_bits_addr_block = GEN_19;
  assign GEN_1_bits_client_xact_id = GEN_20;
  assign GEN_1_bits_addr_beat = GEN_21;
  assign GEN_1_bits_is_builtin_type = GEN_22;
  assign GEN_1_bits_a_type = GEN_23;
  assign GEN_1_bits_union = GEN_24;
  assign GEN_1_bits_data = GEN_25;
  assign GEN_2_ready = GEN_17;
  assign GEN_2_valid = GEN_18;
  assign GEN_2_bits_addr_block = GEN_19;
  assign GEN_2_bits_client_xact_id = GEN_20;
  assign GEN_2_bits_addr_beat = GEN_21;
  assign GEN_2_bits_is_builtin_type = GEN_22;
  assign GEN_2_bits_a_type = GEN_23;
  assign GEN_2_bits_union = GEN_24;
  assign GEN_2_bits_data = GEN_25;
  assign GEN_3_ready = GEN_17;
  assign GEN_3_valid = GEN_18;
  assign GEN_3_bits_addr_block = GEN_19;
  assign GEN_3_bits_client_xact_id = GEN_20;
  assign GEN_3_bits_addr_beat = GEN_21;
  assign GEN_3_bits_is_builtin_type = GEN_22;
  assign GEN_3_bits_a_type = GEN_23;
  assign GEN_3_bits_union = GEN_24;
  assign GEN_3_bits_data = GEN_25;
  assign GEN_4_ready = GEN_17;
  assign GEN_4_valid = GEN_18;
  assign GEN_4_bits_addr_block = GEN_19;
  assign GEN_4_bits_client_xact_id = GEN_20;
  assign GEN_4_bits_addr_beat = GEN_21;
  assign GEN_4_bits_is_builtin_type = GEN_22;
  assign GEN_4_bits_a_type = GEN_23;
  assign GEN_4_bits_union = GEN_24;
  assign GEN_4_bits_data = GEN_25;
  assign GEN_5_ready = GEN_17;
  assign GEN_5_valid = GEN_18;
  assign GEN_5_bits_addr_block = GEN_19;
  assign GEN_5_bits_client_xact_id = GEN_20;
  assign GEN_5_bits_addr_beat = GEN_21;
  assign GEN_5_bits_is_builtin_type = GEN_22;
  assign GEN_5_bits_a_type = GEN_23;
  assign GEN_5_bits_union = GEN_24;
  assign GEN_5_bits_data = GEN_25;
  assign GEN_6_ready = GEN_17;
  assign GEN_6_valid = GEN_18;
  assign GEN_6_bits_addr_block = GEN_19;
  assign GEN_6_bits_client_xact_id = GEN_20;
  assign GEN_6_bits_addr_beat = GEN_21;
  assign GEN_6_bits_is_builtin_type = GEN_22;
  assign GEN_6_bits_a_type = GEN_23;
  assign GEN_6_bits_union = GEN_24;
  assign GEN_6_bits_data = GEN_25;
  assign GEN_7_ready = GEN_17;
  assign GEN_7_valid = GEN_18;
  assign GEN_7_bits_addr_block = GEN_19;
  assign GEN_7_bits_client_xact_id = GEN_20;
  assign GEN_7_bits_addr_beat = GEN_21;
  assign GEN_7_bits_is_builtin_type = GEN_22;
  assign GEN_7_bits_a_type = GEN_23;
  assign GEN_7_bits_union = GEN_24;
  assign GEN_7_bits_data = GEN_25;
  assign T_886 = T_882 != 3'h0;
  assign T_895_0 = 3'h3;
  assign T_897 = io_out_bits_a_type == T_895_0;
  assign T_898 = io_out_bits_is_builtin_type & T_897;
  assign T_899 = io_out_ready & io_out_valid;
  assign T_900 = T_899 & T_898;
  assign T_904 = T_882 + 3'h1;
  assign T_905 = T_904[2:0];
  assign GEN_152 = T_900 ? io_chosen : T_884;
  assign GEN_153 = T_900 ? T_905 : T_882;
  assign GEN_154 = T_886 ? T_884 : choice;
  assign GEN_155 = T_899 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign T_912 = validMask_1 | validMask_2;
  assign T_913 = T_912 | io_in_0_valid;
  assign T_914 = T_913 | io_in_1_valid;
  assign T_918 = validMask_1 == 1'h0;
  assign T_920 = T_912 == 1'h0;
  assign T_922 = T_913 == 1'h0;
  assign T_924 = T_914 == 1'h0;
  assign T_928 = grantMask_1 | T_922;
  assign T_929 = T_918 & grantMask_2;
  assign T_930 = T_929 | T_924;
  assign T_932 = T_884 == 2'h0;
  assign T_933 = T_886 ? T_932 : T_920;
  assign T_934 = T_933 & io_out_ready;
  assign T_936 = T_884 == 2'h1;
  assign T_937 = T_886 ? T_936 : T_928;
  assign T_938 = T_937 & io_out_ready;
  assign T_940 = T_884 == 2'h2;
  assign T_941 = T_886 ? T_940 : T_930;
  assign T_942 = T_941 & io_out_ready;
  assign GEN_156 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_157 = io_in_0_valid ? 2'h0 : GEN_156;
  assign GEN_158 = validMask_2 ? 2'h2 : GEN_157;
  assign GEN_159 = validMask_1 ? 2'h1 : GEN_158;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_882 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_884 = GEN_1[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_882 <= 3'h0;
    end else begin
      if(T_900) begin
        T_882 <= T_905;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_900) begin
        T_884 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_899) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module LockingRRArbiter_6(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_voluntary,
  input  [2:0] io_in_0_bits_r_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_voluntary,
  input  [2:0] io_in_1_bits_r_type,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [25:0] io_in_2_bits_addr_block,
  input  [1:0] io_in_2_bits_client_xact_id,
  input   io_in_2_bits_voluntary,
  input  [2:0] io_in_2_bits_r_type,
  input  [63:0] io_in_2_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_voluntary,
  output [2:0] io_out_bits_r_type,
  output [63:0] io_out_bits_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [25:0] GEN_0_bits_addr_block;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire  GEN_0_bits_voluntary;
  wire [2:0] GEN_0_bits_r_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [25:0] GEN_10;
  wire [1:0] GEN_11;
  wire  GEN_12;
  wire [2:0] GEN_13;
  wire [63:0] GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [25:0] GEN_18;
  wire [1:0] GEN_19;
  wire  GEN_20;
  wire [2:0] GEN_21;
  wire [63:0] GEN_22;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [25:0] GEN_1_bits_addr_block;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire  GEN_1_bits_voluntary;
  wire [2:0] GEN_1_bits_r_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [25:0] GEN_2_bits_addr_block;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire  GEN_2_bits_voluntary;
  wire [2:0] GEN_2_bits_r_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [25:0] GEN_3_bits_addr_block;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire  GEN_3_bits_voluntary;
  wire [2:0] GEN_3_bits_r_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [25:0] GEN_4_bits_addr_block;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire  GEN_4_bits_voluntary;
  wire [2:0] GEN_4_bits_r_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [25:0] GEN_5_bits_addr_block;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire  GEN_5_bits_voluntary;
  wire [2:0] GEN_5_bits_r_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [25:0] GEN_6_bits_addr_block;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire  GEN_6_bits_voluntary;
  wire [2:0] GEN_6_bits_r_type;
  wire [63:0] GEN_6_bits_data;
  reg [2:0] T_852;
  reg [31:0] GEN_0;
  reg [1:0] T_854;
  reg [31:0] GEN_1;
  wire  T_856;
  wire  T_858;
  wire  T_859;
  wire  T_860;
  wire  T_861;
  wire  T_862;
  wire  T_864;
  wire  T_865;
  wire [3:0] T_869;
  wire [2:0] T_870;
  wire [1:0] GEN_119;
  wire [2:0] GEN_120;
  wire [1:0] GEN_121;
  reg [1:0] lastGrant;
  reg [31:0] GEN_2;
  wire [1:0] GEN_122;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  validMask_1;
  wire  validMask_2;
  wire  T_877;
  wire  T_878;
  wire  T_879;
  wire  T_883;
  wire  T_885;
  wire  T_887;
  wire  T_889;
  wire  T_893;
  wire  T_894;
  wire  T_895;
  wire  T_897;
  wire  T_898;
  wire  T_899;
  wire  T_901;
  wire  T_902;
  wire  T_903;
  wire  T_905;
  wire  T_906;
  wire  T_907;
  wire [1:0] GEN_123;
  wire [1:0] GEN_124;
  wire [1:0] GEN_125;
  wire [1:0] GEN_126;
  assign io_in_0_ready = T_899;
  assign io_in_1_ready = T_903;
  assign io_in_2_ready = T_907;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_addr_block = GEN_2_bits_addr_block;
  assign io_out_bits_client_xact_id = GEN_3_bits_client_xact_id;
  assign io_out_bits_voluntary = GEN_4_bits_voluntary;
  assign io_out_bits_r_type = GEN_5_bits_r_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_chosen = GEN_121;
  assign choice = GEN_126;
  assign GEN_0_ready = GEN_15;
  assign GEN_0_valid = GEN_16;
  assign GEN_0_bits_addr_beat = GEN_17;
  assign GEN_0_bits_addr_block = GEN_18;
  assign GEN_0_bits_client_xact_id = GEN_19;
  assign GEN_0_bits_voluntary = GEN_20;
  assign GEN_0_bits_r_type = GEN_21;
  assign GEN_0_bits_data = GEN_22;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_15 = 2'h2 == io_chosen ? io_in_2_ready : GEN_7;
  assign GEN_16 = 2'h2 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_9;
  assign GEN_18 = 2'h2 == io_chosen ? io_in_2_bits_addr_block : GEN_10;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_11;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_voluntary : GEN_12;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_r_type : GEN_13;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_data : GEN_14;
  assign GEN_1_ready = GEN_15;
  assign GEN_1_valid = GEN_16;
  assign GEN_1_bits_addr_beat = GEN_17;
  assign GEN_1_bits_addr_block = GEN_18;
  assign GEN_1_bits_client_xact_id = GEN_19;
  assign GEN_1_bits_voluntary = GEN_20;
  assign GEN_1_bits_r_type = GEN_21;
  assign GEN_1_bits_data = GEN_22;
  assign GEN_2_ready = GEN_15;
  assign GEN_2_valid = GEN_16;
  assign GEN_2_bits_addr_beat = GEN_17;
  assign GEN_2_bits_addr_block = GEN_18;
  assign GEN_2_bits_client_xact_id = GEN_19;
  assign GEN_2_bits_voluntary = GEN_20;
  assign GEN_2_bits_r_type = GEN_21;
  assign GEN_2_bits_data = GEN_22;
  assign GEN_3_ready = GEN_15;
  assign GEN_3_valid = GEN_16;
  assign GEN_3_bits_addr_beat = GEN_17;
  assign GEN_3_bits_addr_block = GEN_18;
  assign GEN_3_bits_client_xact_id = GEN_19;
  assign GEN_3_bits_voluntary = GEN_20;
  assign GEN_3_bits_r_type = GEN_21;
  assign GEN_3_bits_data = GEN_22;
  assign GEN_4_ready = GEN_15;
  assign GEN_4_valid = GEN_16;
  assign GEN_4_bits_addr_beat = GEN_17;
  assign GEN_4_bits_addr_block = GEN_18;
  assign GEN_4_bits_client_xact_id = GEN_19;
  assign GEN_4_bits_voluntary = GEN_20;
  assign GEN_4_bits_r_type = GEN_21;
  assign GEN_4_bits_data = GEN_22;
  assign GEN_5_ready = GEN_15;
  assign GEN_5_valid = GEN_16;
  assign GEN_5_bits_addr_beat = GEN_17;
  assign GEN_5_bits_addr_block = GEN_18;
  assign GEN_5_bits_client_xact_id = GEN_19;
  assign GEN_5_bits_voluntary = GEN_20;
  assign GEN_5_bits_r_type = GEN_21;
  assign GEN_5_bits_data = GEN_22;
  assign GEN_6_ready = GEN_15;
  assign GEN_6_valid = GEN_16;
  assign GEN_6_bits_addr_beat = GEN_17;
  assign GEN_6_bits_addr_block = GEN_18;
  assign GEN_6_bits_client_xact_id = GEN_19;
  assign GEN_6_bits_voluntary = GEN_20;
  assign GEN_6_bits_r_type = GEN_21;
  assign GEN_6_bits_data = GEN_22;
  assign T_856 = T_852 != 3'h0;
  assign T_858 = io_out_bits_r_type == 3'h0;
  assign T_859 = io_out_bits_r_type == 3'h1;
  assign T_860 = io_out_bits_r_type == 3'h2;
  assign T_861 = T_858 | T_859;
  assign T_862 = T_861 | T_860;
  assign T_864 = io_out_ready & io_out_valid;
  assign T_865 = T_864 & T_862;
  assign T_869 = T_852 + 3'h1;
  assign T_870 = T_869[2:0];
  assign GEN_119 = T_865 ? io_chosen : T_854;
  assign GEN_120 = T_865 ? T_870 : T_852;
  assign GEN_121 = T_856 ? T_854 : choice;
  assign GEN_122 = T_864 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign T_877 = validMask_1 | validMask_2;
  assign T_878 = T_877 | io_in_0_valid;
  assign T_879 = T_878 | io_in_1_valid;
  assign T_883 = validMask_1 == 1'h0;
  assign T_885 = T_877 == 1'h0;
  assign T_887 = T_878 == 1'h0;
  assign T_889 = T_879 == 1'h0;
  assign T_893 = grantMask_1 | T_887;
  assign T_894 = T_883 & grantMask_2;
  assign T_895 = T_894 | T_889;
  assign T_897 = T_854 == 2'h0;
  assign T_898 = T_856 ? T_897 : T_885;
  assign T_899 = T_898 & io_out_ready;
  assign T_901 = T_854 == 2'h1;
  assign T_902 = T_856 ? T_901 : T_893;
  assign T_903 = T_902 & io_out_ready;
  assign T_905 = T_854 == 2'h2;
  assign T_906 = T_856 ? T_905 : T_895;
  assign T_907 = T_906 & io_out_ready;
  assign GEN_123 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_124 = io_in_0_valid ? 2'h0 : GEN_123;
  assign GEN_125 = validMask_2 ? 2'h2 : GEN_124;
  assign GEN_126 = validMask_1 ? 2'h1 : GEN_125;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_852 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_854 = GEN_1[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_852 <= 3'h0;
    end else begin
      if(T_865) begin
        T_852 <= T_870;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_865) begin
        T_854 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_864) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientTileLinkIOArbiter(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_probe_ready,
  output  io_in_0_probe_valid,
  output [25:0] io_in_0_probe_bits_addr_block,
  output [1:0] io_in_0_probe_bits_p_type,
  output  io_in_0_release_ready,
  input   io_in_0_release_valid,
  input  [2:0] io_in_0_release_bits_addr_beat,
  input  [25:0] io_in_0_release_bits_addr_block,
  input  [1:0] io_in_0_release_bits_client_xact_id,
  input   io_in_0_release_bits_voluntary,
  input  [2:0] io_in_0_release_bits_r_type,
  input  [63:0] io_in_0_release_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  output  io_in_0_grant_bits_manager_id,
  output  io_in_0_finish_ready,
  input   io_in_0_finish_valid,
  input   io_in_0_finish_bits_manager_xact_id,
  input   io_in_0_finish_bits_manager_id,
  output  io_in_1_acquire_ready,
  input   io_in_1_acquire_valid,
  input  [25:0] io_in_1_acquire_bits_addr_block,
  input  [1:0] io_in_1_acquire_bits_client_xact_id,
  input  [2:0] io_in_1_acquire_bits_addr_beat,
  input   io_in_1_acquire_bits_is_builtin_type,
  input  [2:0] io_in_1_acquire_bits_a_type,
  input  [10:0] io_in_1_acquire_bits_union,
  input  [63:0] io_in_1_acquire_bits_data,
  input   io_in_1_probe_ready,
  output  io_in_1_probe_valid,
  output [25:0] io_in_1_probe_bits_addr_block,
  output [1:0] io_in_1_probe_bits_p_type,
  output  io_in_1_release_ready,
  input   io_in_1_release_valid,
  input  [2:0] io_in_1_release_bits_addr_beat,
  input  [25:0] io_in_1_release_bits_addr_block,
  input  [1:0] io_in_1_release_bits_client_xact_id,
  input   io_in_1_release_bits_voluntary,
  input  [2:0] io_in_1_release_bits_r_type,
  input  [63:0] io_in_1_release_bits_data,
  input   io_in_1_grant_ready,
  output  io_in_1_grant_valid,
  output [2:0] io_in_1_grant_bits_addr_beat,
  output [1:0] io_in_1_grant_bits_client_xact_id,
  output  io_in_1_grant_bits_manager_xact_id,
  output  io_in_1_grant_bits_is_builtin_type,
  output [3:0] io_in_1_grant_bits_g_type,
  output [63:0] io_in_1_grant_bits_data,
  output  io_in_1_grant_bits_manager_id,
  output  io_in_1_finish_ready,
  input   io_in_1_finish_valid,
  input   io_in_1_finish_bits_manager_xact_id,
  input   io_in_1_finish_bits_manager_id,
  output  io_in_2_acquire_ready,
  input   io_in_2_acquire_valid,
  input  [25:0] io_in_2_acquire_bits_addr_block,
  input  [1:0] io_in_2_acquire_bits_client_xact_id,
  input  [2:0] io_in_2_acquire_bits_addr_beat,
  input   io_in_2_acquire_bits_is_builtin_type,
  input  [2:0] io_in_2_acquire_bits_a_type,
  input  [10:0] io_in_2_acquire_bits_union,
  input  [63:0] io_in_2_acquire_bits_data,
  input   io_in_2_probe_ready,
  output  io_in_2_probe_valid,
  output [25:0] io_in_2_probe_bits_addr_block,
  output [1:0] io_in_2_probe_bits_p_type,
  output  io_in_2_release_ready,
  input   io_in_2_release_valid,
  input  [2:0] io_in_2_release_bits_addr_beat,
  input  [25:0] io_in_2_release_bits_addr_block,
  input  [1:0] io_in_2_release_bits_client_xact_id,
  input   io_in_2_release_bits_voluntary,
  input  [2:0] io_in_2_release_bits_r_type,
  input  [63:0] io_in_2_release_bits_data,
  input   io_in_2_grant_ready,
  output  io_in_2_grant_valid,
  output [2:0] io_in_2_grant_bits_addr_beat,
  output [1:0] io_in_2_grant_bits_client_xact_id,
  output  io_in_2_grant_bits_manager_xact_id,
  output  io_in_2_grant_bits_is_builtin_type,
  output [3:0] io_in_2_grant_bits_g_type,
  output [63:0] io_in_2_grant_bits_data,
  output  io_in_2_grant_bits_manager_id,
  output  io_in_2_finish_ready,
  input   io_in_2_finish_valid,
  input   io_in_2_finish_bits_manager_xact_id,
  input   io_in_2_finish_bits_manager_id,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [1:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [10:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_probe_ready,
  input   io_out_probe_valid,
  input  [25:0] io_out_probe_bits_addr_block,
  input  [1:0] io_out_probe_bits_p_type,
  input   io_out_release_ready,
  output  io_out_release_valid,
  output [2:0] io_out_release_bits_addr_beat,
  output [25:0] io_out_release_bits_addr_block,
  output [1:0] io_out_release_bits_client_xact_id,
  output  io_out_release_bits_voluntary,
  output [2:0] io_out_release_bits_r_type,
  output [63:0] io_out_release_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [1:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data,
  input   io_out_grant_bits_manager_id,
  input   io_out_finish_ready,
  output  io_out_finish_valid,
  output  io_out_finish_bits_manager_xact_id,
  output  io_out_finish_bits_manager_id
);
  wire  LockingRRArbiter_5_1_clk;
  wire  LockingRRArbiter_5_1_reset;
  wire  LockingRRArbiter_5_1_io_in_0_ready;
  wire  LockingRRArbiter_5_1_io_in_0_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_0_bits_addr_block;
  wire [1:0] LockingRRArbiter_5_1_io_in_0_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_0_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_0_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_0_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_in_0_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_0_bits_data;
  wire  LockingRRArbiter_5_1_io_in_1_ready;
  wire  LockingRRArbiter_5_1_io_in_1_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_1_bits_addr_block;
  wire [1:0] LockingRRArbiter_5_1_io_in_1_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_1_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_1_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_1_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_in_1_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_1_bits_data;
  wire  LockingRRArbiter_5_1_io_in_2_ready;
  wire  LockingRRArbiter_5_1_io_in_2_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_2_bits_addr_block;
  wire [1:0] LockingRRArbiter_5_1_io_in_2_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_2_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_2_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_2_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_in_2_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_2_bits_data;
  wire  LockingRRArbiter_5_1_io_out_ready;
  wire  LockingRRArbiter_5_1_io_out_valid;
  wire [25:0] LockingRRArbiter_5_1_io_out_bits_addr_block;
  wire [1:0] LockingRRArbiter_5_1_io_out_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_out_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_out_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_out_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_out_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_out_bits_data;
  wire [1:0] LockingRRArbiter_5_1_io_chosen;
  wire [3:0] T_6920;
  wire [3:0] T_6922;
  wire [3:0] T_6924;
  wire  LockingRRArbiter_6_1_clk;
  wire  LockingRRArbiter_6_1_reset;
  wire  LockingRRArbiter_6_1_io_in_0_ready;
  wire  LockingRRArbiter_6_1_io_in_0_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_0_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_0_bits_addr_block;
  wire [1:0] LockingRRArbiter_6_1_io_in_0_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_0_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_0_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_0_bits_data;
  wire  LockingRRArbiter_6_1_io_in_1_ready;
  wire  LockingRRArbiter_6_1_io_in_1_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_1_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_1_bits_addr_block;
  wire [1:0] LockingRRArbiter_6_1_io_in_1_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_1_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_1_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_1_bits_data;
  wire  LockingRRArbiter_6_1_io_in_2_ready;
  wire  LockingRRArbiter_6_1_io_in_2_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_2_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_2_bits_addr_block;
  wire [1:0] LockingRRArbiter_6_1_io_in_2_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_2_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_2_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_2_bits_data;
  wire  LockingRRArbiter_6_1_io_out_ready;
  wire  LockingRRArbiter_6_1_io_out_valid;
  wire [2:0] LockingRRArbiter_6_1_io_out_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_out_bits_addr_block;
  wire [1:0] LockingRRArbiter_6_1_io_out_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_out_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_out_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_out_bits_data;
  wire [1:0] LockingRRArbiter_6_1_io_chosen;
  wire [3:0] T_6926;
  wire [3:0] T_6928;
  wire [3:0] T_6930;
  wire  T_6931;
  wire  T_6932;
  wire  T_6937;
  wire  GEN_0;
  wire  GEN_1;
  wire  T_6942;
  wire  GEN_2;
  wire  GEN_3;
  wire  T_6947;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  reg [31:0] GEN_12;
  wire  GEN_7;
  reg [31:0] GEN_13;
  wire  GEN_8;
  reg [31:0] GEN_14;
  wire  GEN_9;
  reg [31:0] GEN_15;
  wire  GEN_10;
  reg [31:0] GEN_16;
  wire  GEN_11;
  reg [31:0] GEN_17;
  LockingRRArbiter_5 LockingRRArbiter_5_1 (
    .clk(LockingRRArbiter_5_1_clk),
    .reset(LockingRRArbiter_5_1_reset),
    .io_in_0_ready(LockingRRArbiter_5_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_5_1_io_in_0_valid),
    .io_in_0_bits_addr_block(LockingRRArbiter_5_1_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_5_1_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(LockingRRArbiter_5_1_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(LockingRRArbiter_5_1_io_in_0_bits_a_type),
    .io_in_0_bits_union(LockingRRArbiter_5_1_io_in_0_bits_union),
    .io_in_0_bits_data(LockingRRArbiter_5_1_io_in_0_bits_data),
    .io_in_1_ready(LockingRRArbiter_5_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_5_1_io_in_1_valid),
    .io_in_1_bits_addr_block(LockingRRArbiter_5_1_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_5_1_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(LockingRRArbiter_5_1_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(LockingRRArbiter_5_1_io_in_1_bits_a_type),
    .io_in_1_bits_union(LockingRRArbiter_5_1_io_in_1_bits_union),
    .io_in_1_bits_data(LockingRRArbiter_5_1_io_in_1_bits_data),
    .io_in_2_ready(LockingRRArbiter_5_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_5_1_io_in_2_valid),
    .io_in_2_bits_addr_block(LockingRRArbiter_5_1_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_5_1_io_in_2_bits_client_xact_id),
    .io_in_2_bits_addr_beat(LockingRRArbiter_5_1_io_in_2_bits_addr_beat),
    .io_in_2_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_a_type(LockingRRArbiter_5_1_io_in_2_bits_a_type),
    .io_in_2_bits_union(LockingRRArbiter_5_1_io_in_2_bits_union),
    .io_in_2_bits_data(LockingRRArbiter_5_1_io_in_2_bits_data),
    .io_out_ready(LockingRRArbiter_5_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_5_1_io_out_valid),
    .io_out_bits_addr_block(LockingRRArbiter_5_1_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(LockingRRArbiter_5_1_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(LockingRRArbiter_5_1_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(LockingRRArbiter_5_1_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(LockingRRArbiter_5_1_io_out_bits_a_type),
    .io_out_bits_union(LockingRRArbiter_5_1_io_out_bits_union),
    .io_out_bits_data(LockingRRArbiter_5_1_io_out_bits_data),
    .io_chosen(LockingRRArbiter_5_1_io_chosen)
  );
  LockingRRArbiter_6 LockingRRArbiter_6_1 (
    .clk(LockingRRArbiter_6_1_clk),
    .reset(LockingRRArbiter_6_1_reset),
    .io_in_0_ready(LockingRRArbiter_6_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_6_1_io_in_0_valid),
    .io_in_0_bits_addr_beat(LockingRRArbiter_6_1_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(LockingRRArbiter_6_1_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_6_1_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(LockingRRArbiter_6_1_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(LockingRRArbiter_6_1_io_in_0_bits_r_type),
    .io_in_0_bits_data(LockingRRArbiter_6_1_io_in_0_bits_data),
    .io_in_1_ready(LockingRRArbiter_6_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_6_1_io_in_1_valid),
    .io_in_1_bits_addr_beat(LockingRRArbiter_6_1_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(LockingRRArbiter_6_1_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_6_1_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(LockingRRArbiter_6_1_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(LockingRRArbiter_6_1_io_in_1_bits_r_type),
    .io_in_1_bits_data(LockingRRArbiter_6_1_io_in_1_bits_data),
    .io_in_2_ready(LockingRRArbiter_6_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_6_1_io_in_2_valid),
    .io_in_2_bits_addr_beat(LockingRRArbiter_6_1_io_in_2_bits_addr_beat),
    .io_in_2_bits_addr_block(LockingRRArbiter_6_1_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_6_1_io_in_2_bits_client_xact_id),
    .io_in_2_bits_voluntary(LockingRRArbiter_6_1_io_in_2_bits_voluntary),
    .io_in_2_bits_r_type(LockingRRArbiter_6_1_io_in_2_bits_r_type),
    .io_in_2_bits_data(LockingRRArbiter_6_1_io_in_2_bits_data),
    .io_out_ready(LockingRRArbiter_6_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_6_1_io_out_valid),
    .io_out_bits_addr_beat(LockingRRArbiter_6_1_io_out_bits_addr_beat),
    .io_out_bits_addr_block(LockingRRArbiter_6_1_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(LockingRRArbiter_6_1_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(LockingRRArbiter_6_1_io_out_bits_voluntary),
    .io_out_bits_r_type(LockingRRArbiter_6_1_io_out_bits_r_type),
    .io_out_bits_data(LockingRRArbiter_6_1_io_out_bits_data),
    .io_chosen(LockingRRArbiter_6_1_io_chosen)
  );
  assign io_in_0_acquire_ready = LockingRRArbiter_5_1_io_in_0_ready;
  assign io_in_0_probe_valid = io_out_probe_valid;
  assign io_in_0_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_0_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_0_release_ready = LockingRRArbiter_6_1_io_in_0_ready;
  assign io_in_0_grant_valid = GEN_0;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = 2'h0;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_in_0_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_0_finish_ready = GEN_6;
  assign io_in_1_acquire_ready = LockingRRArbiter_5_1_io_in_1_ready;
  assign io_in_1_probe_valid = io_out_probe_valid;
  assign io_in_1_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_1_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_1_release_ready = LockingRRArbiter_6_1_io_in_1_ready;
  assign io_in_1_grant_valid = GEN_2;
  assign io_in_1_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_1_grant_bits_client_xact_id = 2'h0;
  assign io_in_1_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_1_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_1_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_1_grant_bits_data = io_out_grant_bits_data;
  assign io_in_1_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_1_finish_ready = GEN_7;
  assign io_in_2_acquire_ready = LockingRRArbiter_5_1_io_in_2_ready;
  assign io_in_2_probe_valid = io_out_probe_valid;
  assign io_in_2_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_2_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_2_release_ready = LockingRRArbiter_6_1_io_in_2_ready;
  assign io_in_2_grant_valid = GEN_4;
  assign io_in_2_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_2_grant_bits_client_xact_id = 2'h0;
  assign io_in_2_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_2_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_2_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_2_grant_bits_data = io_out_grant_bits_data;
  assign io_in_2_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_2_finish_ready = GEN_8;
  assign io_out_acquire_valid = LockingRRArbiter_5_1_io_out_valid;
  assign io_out_acquire_bits_addr_block = LockingRRArbiter_5_1_io_out_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = LockingRRArbiter_5_1_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = LockingRRArbiter_5_1_io_out_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = LockingRRArbiter_5_1_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = LockingRRArbiter_5_1_io_out_bits_a_type;
  assign io_out_acquire_bits_union = LockingRRArbiter_5_1_io_out_bits_union;
  assign io_out_acquire_bits_data = LockingRRArbiter_5_1_io_out_bits_data;
  assign io_out_probe_ready = T_6932;
  assign io_out_release_valid = LockingRRArbiter_6_1_io_out_valid;
  assign io_out_release_bits_addr_beat = LockingRRArbiter_6_1_io_out_bits_addr_beat;
  assign io_out_release_bits_addr_block = LockingRRArbiter_6_1_io_out_bits_addr_block;
  assign io_out_release_bits_client_xact_id = LockingRRArbiter_6_1_io_out_bits_client_xact_id;
  assign io_out_release_bits_voluntary = LockingRRArbiter_6_1_io_out_bits_voluntary;
  assign io_out_release_bits_r_type = LockingRRArbiter_6_1_io_out_bits_r_type;
  assign io_out_release_bits_data = LockingRRArbiter_6_1_io_out_bits_data;
  assign io_out_grant_ready = GEN_5;
  assign io_out_finish_valid = GEN_9;
  assign io_out_finish_bits_manager_xact_id = GEN_10;
  assign io_out_finish_bits_manager_id = GEN_11;
  assign LockingRRArbiter_5_1_clk = clk;
  assign LockingRRArbiter_5_1_reset = reset;
  assign LockingRRArbiter_5_1_io_in_0_valid = io_in_0_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_0_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_0_bits_client_xact_id = T_6920[1:0];
  assign LockingRRArbiter_5_1_io_in_0_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_0_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_0_bits_a_type = io_in_0_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_0_bits_union = io_in_0_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_0_bits_data = io_in_0_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_1_valid = io_in_1_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_1_bits_addr_block = io_in_1_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_1_bits_client_xact_id = T_6922[1:0];
  assign LockingRRArbiter_5_1_io_in_1_bits_addr_beat = io_in_1_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_1_bits_is_builtin_type = io_in_1_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_1_bits_a_type = io_in_1_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_1_bits_union = io_in_1_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_1_bits_data = io_in_1_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_2_valid = io_in_2_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_2_bits_addr_block = io_in_2_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_2_bits_client_xact_id = T_6924[1:0];
  assign LockingRRArbiter_5_1_io_in_2_bits_addr_beat = io_in_2_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_2_bits_is_builtin_type = io_in_2_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_2_bits_a_type = io_in_2_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_2_bits_union = io_in_2_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_2_bits_data = io_in_2_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_out_ready = io_out_acquire_ready;
  assign T_6920 = {io_in_0_acquire_bits_client_xact_id,2'h0};
  assign T_6922 = {io_in_1_acquire_bits_client_xact_id,2'h1};
  assign T_6924 = {io_in_2_acquire_bits_client_xact_id,2'h2};
  assign LockingRRArbiter_6_1_clk = clk;
  assign LockingRRArbiter_6_1_reset = reset;
  assign LockingRRArbiter_6_1_io_in_0_valid = io_in_0_release_valid;
  assign LockingRRArbiter_6_1_io_in_0_bits_addr_beat = io_in_0_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_0_bits_addr_block = io_in_0_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_0_bits_client_xact_id = T_6926[1:0];
  assign LockingRRArbiter_6_1_io_in_0_bits_voluntary = io_in_0_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_0_bits_r_type = io_in_0_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_0_bits_data = io_in_0_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_1_valid = io_in_1_release_valid;
  assign LockingRRArbiter_6_1_io_in_1_bits_addr_beat = io_in_1_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_1_bits_addr_block = io_in_1_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_1_bits_client_xact_id = T_6928[1:0];
  assign LockingRRArbiter_6_1_io_in_1_bits_voluntary = io_in_1_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_1_bits_r_type = io_in_1_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_1_bits_data = io_in_1_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_2_valid = io_in_2_release_valid;
  assign LockingRRArbiter_6_1_io_in_2_bits_addr_beat = io_in_2_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_2_bits_addr_block = io_in_2_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_2_bits_client_xact_id = T_6930[1:0];
  assign LockingRRArbiter_6_1_io_in_2_bits_voluntary = io_in_2_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_2_bits_r_type = io_in_2_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_2_bits_data = io_in_2_release_bits_data;
  assign LockingRRArbiter_6_1_io_out_ready = io_out_release_ready;
  assign T_6926 = {io_in_0_release_bits_client_xact_id,2'h0};
  assign T_6928 = {io_in_1_release_bits_client_xact_id,2'h1};
  assign T_6930 = {io_in_2_release_bits_client_xact_id,2'h2};
  assign T_6931 = io_in_0_probe_ready & io_in_1_probe_ready;
  assign T_6932 = T_6931 & io_in_2_probe_ready;
  assign T_6937 = io_out_grant_bits_client_xact_id == 2'h0;
  assign GEN_0 = T_6937 ? io_out_grant_valid : 1'h0;
  assign GEN_1 = T_6937 ? io_in_0_grant_ready : 1'h0;
  assign T_6942 = io_out_grant_bits_client_xact_id == 2'h1;
  assign GEN_2 = T_6942 ? io_out_grant_valid : 1'h0;
  assign GEN_3 = T_6942 ? io_in_1_grant_ready : GEN_1;
  assign T_6947 = io_out_grant_bits_client_xact_id == 2'h2;
  assign GEN_4 = T_6947 ? io_out_grant_valid : 1'h0;
  assign GEN_5 = T_6947 ? io_in_2_grant_ready : GEN_3;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_6 = GEN_12[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_7 = GEN_13[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_8 = GEN_14[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_9 = GEN_15[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_10 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_11 = GEN_17[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_12 = {1{$random}};
  GEN_13 = {1{$random}};
  GEN_14 = {1{$random}};
  GEN_15 = {1{$random}};
  GEN_16 = {1{$random}};
  GEN_17 = {1{$random}};
  end
`endif
endmodule
module LockingRRArbiter_7(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_p_type,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_p_type,
  input   io_in_1_bits_client_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [1:0] io_in_2_bits_p_type,
  input   io_in_2_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_p_type,
  output  io_out_bits_client_id,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [25:0] GEN_0_bits_addr_block;
  wire [1:0] GEN_0_bits_p_type;
  wire  GEN_0_bits_client_id;
  wire  GEN_4;
  wire  GEN_5;
  wire [25:0] GEN_6;
  wire [1:0] GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [25:0] GEN_11;
  wire [1:0] GEN_12;
  wire  GEN_13;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [25:0] GEN_1_bits_addr_block;
  wire [1:0] GEN_1_bits_p_type;
  wire  GEN_1_bits_client_id;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [25:0] GEN_2_bits_addr_block;
  wire [1:0] GEN_2_bits_p_type;
  wire  GEN_2_bits_client_id;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [25:0] GEN_3_bits_addr_block;
  wire [1:0] GEN_3_bits_p_type;
  wire  GEN_3_bits_client_id;
  reg [2:0] T_762;
  reg [31:0] GEN_0;
  reg [1:0] T_764;
  reg [31:0] GEN_1;
  wire  T_766;
  wire  T_768;
  wire [1:0] GEN_46;
  reg [1:0] lastGrant;
  reg [31:0] GEN_2;
  wire [1:0] GEN_47;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  validMask_1;
  wire  validMask_2;
  wire  T_781;
  wire  T_782;
  wire  T_783;
  wire  T_787;
  wire  T_789;
  wire  T_791;
  wire  T_793;
  wire  T_797;
  wire  T_798;
  wire  T_799;
  wire  T_801;
  wire  T_802;
  wire  T_803;
  wire  T_805;
  wire  T_806;
  wire  T_807;
  wire  T_809;
  wire  T_810;
  wire  T_811;
  wire [1:0] GEN_48;
  wire [1:0] GEN_49;
  wire [1:0] GEN_50;
  wire [1:0] GEN_51;
  assign io_in_0_ready = T_803;
  assign io_in_1_ready = T_807;
  assign io_in_2_ready = T_811;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_block = GEN_1_bits_addr_block;
  assign io_out_bits_p_type = GEN_2_bits_p_type;
  assign io_out_bits_client_id = GEN_3_bits_client_id;
  assign io_chosen = GEN_46;
  assign choice = GEN_51;
  assign GEN_0_ready = GEN_9;
  assign GEN_0_valid = GEN_10;
  assign GEN_0_bits_addr_block = GEN_11;
  assign GEN_0_bits_p_type = GEN_12;
  assign GEN_0_bits_client_id = GEN_13;
  assign GEN_4 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_5 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_6 = 2'h1 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_bits_p_type : io_in_0_bits_p_type;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_9 = 2'h2 == io_chosen ? io_in_2_ready : GEN_4;
  assign GEN_10 = 2'h2 == io_chosen ? io_in_2_valid : GEN_5;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_bits_addr_block : GEN_6;
  assign GEN_12 = 2'h2 == io_chosen ? io_in_2_bits_p_type : GEN_7;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_client_id : GEN_8;
  assign GEN_1_ready = GEN_9;
  assign GEN_1_valid = GEN_10;
  assign GEN_1_bits_addr_block = GEN_11;
  assign GEN_1_bits_p_type = GEN_12;
  assign GEN_1_bits_client_id = GEN_13;
  assign GEN_2_ready = GEN_9;
  assign GEN_2_valid = GEN_10;
  assign GEN_2_bits_addr_block = GEN_11;
  assign GEN_2_bits_p_type = GEN_12;
  assign GEN_2_bits_client_id = GEN_13;
  assign GEN_3_ready = GEN_9;
  assign GEN_3_valid = GEN_10;
  assign GEN_3_bits_addr_block = GEN_11;
  assign GEN_3_bits_p_type = GEN_12;
  assign GEN_3_bits_client_id = GEN_13;
  assign T_766 = T_762 != 3'h0;
  assign T_768 = io_out_ready & io_out_valid;
  assign GEN_46 = T_766 ? T_764 : choice;
  assign GEN_47 = T_768 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign T_781 = validMask_1 | validMask_2;
  assign T_782 = T_781 | io_in_0_valid;
  assign T_783 = T_782 | io_in_1_valid;
  assign T_787 = validMask_1 == 1'h0;
  assign T_789 = T_781 == 1'h0;
  assign T_791 = T_782 == 1'h0;
  assign T_793 = T_783 == 1'h0;
  assign T_797 = grantMask_1 | T_791;
  assign T_798 = T_787 & grantMask_2;
  assign T_799 = T_798 | T_793;
  assign T_801 = T_764 == 2'h0;
  assign T_802 = T_766 ? T_801 : T_789;
  assign T_803 = T_802 & io_out_ready;
  assign T_805 = T_764 == 2'h1;
  assign T_806 = T_766 ? T_805 : T_797;
  assign T_807 = T_806 & io_out_ready;
  assign T_809 = T_764 == 2'h2;
  assign T_810 = T_766 ? T_809 : T_799;
  assign T_811 = T_810 & io_out_ready;
  assign GEN_48 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_49 = io_in_0_valid ? 2'h0 : GEN_48;
  assign GEN_50 = validMask_2 ? 2'h2 : GEN_49;
  assign GEN_51 = validMask_1 ? 2'h1 : GEN_50;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_762 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_764 = GEN_1[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_762 <= 3'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(T_768) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module LockingRRArbiter_8(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_client_xact_id,
  input  [1:0] io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_client_xact_id,
  input  [1:0] io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input   io_in_2_bits_client_xact_id,
  input  [1:0] io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_is_builtin_type,
  input  [3:0] io_in_2_bits_g_type,
  input  [63:0] io_in_2_bits_data,
  input   io_in_2_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_client_xact_id,
  output [1:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire  GEN_0_bits_client_xact_id;
  wire [1:0] GEN_0_bits_manager_xact_id;
  wire  GEN_0_bits_is_builtin_type;
  wire [3:0] GEN_0_bits_g_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_0_bits_client_id;
  wire  GEN_8;
  wire  GEN_9;
  wire [2:0] GEN_10;
  wire  GEN_11;
  wire [1:0] GEN_12;
  wire  GEN_13;
  wire [3:0] GEN_14;
  wire [63:0] GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire  GEN_20;
  wire [1:0] GEN_21;
  wire  GEN_22;
  wire [3:0] GEN_23;
  wire [63:0] GEN_24;
  wire  GEN_25;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire  GEN_1_bits_client_xact_id;
  wire [1:0] GEN_1_bits_manager_xact_id;
  wire  GEN_1_bits_is_builtin_type;
  wire [3:0] GEN_1_bits_g_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_1_bits_client_id;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire  GEN_2_bits_client_xact_id;
  wire [1:0] GEN_2_bits_manager_xact_id;
  wire  GEN_2_bits_is_builtin_type;
  wire [3:0] GEN_2_bits_g_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_2_bits_client_id;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire  GEN_3_bits_client_xact_id;
  wire [1:0] GEN_3_bits_manager_xact_id;
  wire  GEN_3_bits_is_builtin_type;
  wire [3:0] GEN_3_bits_g_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_3_bits_client_id;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire  GEN_4_bits_client_xact_id;
  wire [1:0] GEN_4_bits_manager_xact_id;
  wire  GEN_4_bits_is_builtin_type;
  wire [3:0] GEN_4_bits_g_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_4_bits_client_id;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire  GEN_5_bits_client_xact_id;
  wire [1:0] GEN_5_bits_manager_xact_id;
  wire  GEN_5_bits_is_builtin_type;
  wire [3:0] GEN_5_bits_g_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_5_bits_client_id;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire  GEN_6_bits_client_xact_id;
  wire [1:0] GEN_6_bits_manager_xact_id;
  wire  GEN_6_bits_is_builtin_type;
  wire [3:0] GEN_6_bits_g_type;
  wire [63:0] GEN_6_bits_data;
  wire  GEN_6_bits_client_id;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [2:0] GEN_7_bits_addr_beat;
  wire  GEN_7_bits_client_xact_id;
  wire [1:0] GEN_7_bits_manager_xact_id;
  wire  GEN_7_bits_is_builtin_type;
  wire [3:0] GEN_7_bits_g_type;
  wire [63:0] GEN_7_bits_data;
  wire  GEN_7_bits_client_id;
  reg [2:0] T_882;
  reg [31:0] GEN_1;
  reg [1:0] T_884;
  reg [31:0] GEN_2;
  wire  T_886;
  wire [2:0] T_894_0;
  wire [3:0] GEN_0;
  wire  T_896;
  wire  T_897;
  wire  T_898;
  wire  T_900;
  wire  T_901;
  wire [3:0] T_905;
  wire [2:0] T_906;
  wire [1:0] GEN_152;
  wire [2:0] GEN_153;
  wire [1:0] GEN_154;
  reg [1:0] lastGrant;
  reg [31:0] GEN_3;
  wire [1:0] GEN_155;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  validMask_1;
  wire  validMask_2;
  wire  T_913;
  wire  T_914;
  wire  T_915;
  wire  T_919;
  wire  T_921;
  wire  T_923;
  wire  T_925;
  wire  T_929;
  wire  T_930;
  wire  T_931;
  wire  T_933;
  wire  T_934;
  wire  T_935;
  wire  T_937;
  wire  T_938;
  wire  T_939;
  wire  T_941;
  wire  T_942;
  wire  T_943;
  wire [1:0] GEN_156;
  wire [1:0] GEN_157;
  wire [1:0] GEN_158;
  wire [1:0] GEN_159;
  assign io_in_0_ready = T_935;
  assign io_in_1_ready = T_939;
  assign io_in_2_ready = T_943;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = GEN_3_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_g_type = GEN_5_bits_g_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_out_bits_client_id = GEN_7_bits_client_id;
  assign io_chosen = GEN_154;
  assign choice = GEN_159;
  assign GEN_0_ready = GEN_17;
  assign GEN_0_valid = GEN_18;
  assign GEN_0_bits_addr_beat = GEN_19;
  assign GEN_0_bits_client_xact_id = GEN_20;
  assign GEN_0_bits_manager_xact_id = GEN_21;
  assign GEN_0_bits_is_builtin_type = GEN_22;
  assign GEN_0_bits_g_type = GEN_23;
  assign GEN_0_bits_data = GEN_24;
  assign GEN_0_bits_client_id = GEN_25;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_ready : GEN_8;
  assign GEN_18 = 2'h2 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_10;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_11;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_manager_xact_id : GEN_12;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_13;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_g_type : GEN_14;
  assign GEN_24 = 2'h2 == io_chosen ? io_in_2_bits_data : GEN_15;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_client_id : GEN_16;
  assign GEN_1_ready = GEN_17;
  assign GEN_1_valid = GEN_18;
  assign GEN_1_bits_addr_beat = GEN_19;
  assign GEN_1_bits_client_xact_id = GEN_20;
  assign GEN_1_bits_manager_xact_id = GEN_21;
  assign GEN_1_bits_is_builtin_type = GEN_22;
  assign GEN_1_bits_g_type = GEN_23;
  assign GEN_1_bits_data = GEN_24;
  assign GEN_1_bits_client_id = GEN_25;
  assign GEN_2_ready = GEN_17;
  assign GEN_2_valid = GEN_18;
  assign GEN_2_bits_addr_beat = GEN_19;
  assign GEN_2_bits_client_xact_id = GEN_20;
  assign GEN_2_bits_manager_xact_id = GEN_21;
  assign GEN_2_bits_is_builtin_type = GEN_22;
  assign GEN_2_bits_g_type = GEN_23;
  assign GEN_2_bits_data = GEN_24;
  assign GEN_2_bits_client_id = GEN_25;
  assign GEN_3_ready = GEN_17;
  assign GEN_3_valid = GEN_18;
  assign GEN_3_bits_addr_beat = GEN_19;
  assign GEN_3_bits_client_xact_id = GEN_20;
  assign GEN_3_bits_manager_xact_id = GEN_21;
  assign GEN_3_bits_is_builtin_type = GEN_22;
  assign GEN_3_bits_g_type = GEN_23;
  assign GEN_3_bits_data = GEN_24;
  assign GEN_3_bits_client_id = GEN_25;
  assign GEN_4_ready = GEN_17;
  assign GEN_4_valid = GEN_18;
  assign GEN_4_bits_addr_beat = GEN_19;
  assign GEN_4_bits_client_xact_id = GEN_20;
  assign GEN_4_bits_manager_xact_id = GEN_21;
  assign GEN_4_bits_is_builtin_type = GEN_22;
  assign GEN_4_bits_g_type = GEN_23;
  assign GEN_4_bits_data = GEN_24;
  assign GEN_4_bits_client_id = GEN_25;
  assign GEN_5_ready = GEN_17;
  assign GEN_5_valid = GEN_18;
  assign GEN_5_bits_addr_beat = GEN_19;
  assign GEN_5_bits_client_xact_id = GEN_20;
  assign GEN_5_bits_manager_xact_id = GEN_21;
  assign GEN_5_bits_is_builtin_type = GEN_22;
  assign GEN_5_bits_g_type = GEN_23;
  assign GEN_5_bits_data = GEN_24;
  assign GEN_5_bits_client_id = GEN_25;
  assign GEN_6_ready = GEN_17;
  assign GEN_6_valid = GEN_18;
  assign GEN_6_bits_addr_beat = GEN_19;
  assign GEN_6_bits_client_xact_id = GEN_20;
  assign GEN_6_bits_manager_xact_id = GEN_21;
  assign GEN_6_bits_is_builtin_type = GEN_22;
  assign GEN_6_bits_g_type = GEN_23;
  assign GEN_6_bits_data = GEN_24;
  assign GEN_6_bits_client_id = GEN_25;
  assign GEN_7_ready = GEN_17;
  assign GEN_7_valid = GEN_18;
  assign GEN_7_bits_addr_beat = GEN_19;
  assign GEN_7_bits_client_xact_id = GEN_20;
  assign GEN_7_bits_manager_xact_id = GEN_21;
  assign GEN_7_bits_is_builtin_type = GEN_22;
  assign GEN_7_bits_g_type = GEN_23;
  assign GEN_7_bits_data = GEN_24;
  assign GEN_7_bits_client_id = GEN_25;
  assign T_886 = T_882 != 3'h0;
  assign T_894_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_894_0};
  assign T_896 = io_out_bits_g_type == GEN_0;
  assign T_897 = io_out_bits_g_type == 4'h0;
  assign T_898 = io_out_bits_is_builtin_type ? T_896 : T_897;
  assign T_900 = io_out_ready & io_out_valid;
  assign T_901 = T_900 & T_898;
  assign T_905 = T_882 + 3'h1;
  assign T_906 = T_905[2:0];
  assign GEN_152 = T_901 ? io_chosen : T_884;
  assign GEN_153 = T_901 ? T_906 : T_882;
  assign GEN_154 = T_886 ? T_884 : choice;
  assign GEN_155 = T_900 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign T_913 = validMask_1 | validMask_2;
  assign T_914 = T_913 | io_in_0_valid;
  assign T_915 = T_914 | io_in_1_valid;
  assign T_919 = validMask_1 == 1'h0;
  assign T_921 = T_913 == 1'h0;
  assign T_923 = T_914 == 1'h0;
  assign T_925 = T_915 == 1'h0;
  assign T_929 = grantMask_1 | T_923;
  assign T_930 = T_919 & grantMask_2;
  assign T_931 = T_930 | T_925;
  assign T_933 = T_884 == 2'h0;
  assign T_934 = T_886 ? T_933 : T_921;
  assign T_935 = T_934 & io_out_ready;
  assign T_937 = T_884 == 2'h1;
  assign T_938 = T_886 ? T_937 : T_929;
  assign T_939 = T_938 & io_out_ready;
  assign T_941 = T_884 == 2'h2;
  assign T_942 = T_886 ? T_941 : T_931;
  assign T_943 = T_942 & io_out_ready;
  assign GEN_156 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_157 = io_in_0_valid ? 2'h0 : GEN_156;
  assign GEN_158 = validMask_2 ? 2'h2 : GEN_157;
  assign GEN_159 = validMask_1 ? 2'h1 : GEN_158;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_882 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_884 = GEN_2[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  lastGrant = GEN_3[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_882 <= 3'h0;
    end else begin
      if(T_901) begin
        T_882 <= T_906;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_901) begin
        T_884 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_900) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module L2BroadcastHub(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input   io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output  io_inner_grant_bits_client_xact_id,
  output [1:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [1:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input   io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [1:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id
);
  wire  trackerList_0_clk;
  wire  trackerList_0_reset;
  wire  trackerList_0_io_inner_acquire_ready;
  wire  trackerList_0_io_inner_acquire_valid;
  wire [25:0] trackerList_0_io_inner_acquire_bits_addr_block;
  wire  trackerList_0_io_inner_acquire_bits_client_xact_id;
  wire [2:0] trackerList_0_io_inner_acquire_bits_addr_beat;
  wire  trackerList_0_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_0_io_inner_acquire_bits_a_type;
  wire [10:0] trackerList_0_io_inner_acquire_bits_union;
  wire [63:0] trackerList_0_io_inner_acquire_bits_data;
  wire  trackerList_0_io_inner_acquire_bits_client_id;
  wire  trackerList_0_io_inner_grant_ready;
  wire  trackerList_0_io_inner_grant_valid;
  wire [2:0] trackerList_0_io_inner_grant_bits_addr_beat;
  wire  trackerList_0_io_inner_grant_bits_client_xact_id;
  wire [1:0] trackerList_0_io_inner_grant_bits_manager_xact_id;
  wire  trackerList_0_io_inner_grant_bits_is_builtin_type;
  wire [3:0] trackerList_0_io_inner_grant_bits_g_type;
  wire [63:0] trackerList_0_io_inner_grant_bits_data;
  wire  trackerList_0_io_inner_grant_bits_client_id;
  wire  trackerList_0_io_inner_finish_ready;
  wire  trackerList_0_io_inner_finish_valid;
  wire [1:0] trackerList_0_io_inner_finish_bits_manager_xact_id;
  wire  trackerList_0_io_inner_probe_ready;
  wire  trackerList_0_io_inner_probe_valid;
  wire [25:0] trackerList_0_io_inner_probe_bits_addr_block;
  wire [1:0] trackerList_0_io_inner_probe_bits_p_type;
  wire  trackerList_0_io_inner_probe_bits_client_id;
  wire  trackerList_0_io_inner_release_ready;
  wire  trackerList_0_io_inner_release_valid;
  wire [2:0] trackerList_0_io_inner_release_bits_addr_beat;
  wire [25:0] trackerList_0_io_inner_release_bits_addr_block;
  wire  trackerList_0_io_inner_release_bits_client_xact_id;
  wire  trackerList_0_io_inner_release_bits_voluntary;
  wire [2:0] trackerList_0_io_inner_release_bits_r_type;
  wire [63:0] trackerList_0_io_inner_release_bits_data;
  wire  trackerList_0_io_inner_release_bits_client_id;
  wire  trackerList_0_io_incoherent_0;
  wire  trackerList_0_io_outer_acquire_ready;
  wire  trackerList_0_io_outer_acquire_valid;
  wire [25:0] trackerList_0_io_outer_acquire_bits_addr_block;
  wire [1:0] trackerList_0_io_outer_acquire_bits_client_xact_id;
  wire [2:0] trackerList_0_io_outer_acquire_bits_addr_beat;
  wire  trackerList_0_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_0_io_outer_acquire_bits_a_type;
  wire [10:0] trackerList_0_io_outer_acquire_bits_union;
  wire [63:0] trackerList_0_io_outer_acquire_bits_data;
  wire  trackerList_0_io_outer_probe_ready;
  wire  trackerList_0_io_outer_probe_valid;
  wire [25:0] trackerList_0_io_outer_probe_bits_addr_block;
  wire [1:0] trackerList_0_io_outer_probe_bits_p_type;
  wire  trackerList_0_io_outer_release_ready;
  wire  trackerList_0_io_outer_release_valid;
  wire [2:0] trackerList_0_io_outer_release_bits_addr_beat;
  wire [25:0] trackerList_0_io_outer_release_bits_addr_block;
  wire [1:0] trackerList_0_io_outer_release_bits_client_xact_id;
  wire  trackerList_0_io_outer_release_bits_voluntary;
  wire [2:0] trackerList_0_io_outer_release_bits_r_type;
  wire [63:0] trackerList_0_io_outer_release_bits_data;
  wire  trackerList_0_io_outer_grant_ready;
  wire  trackerList_0_io_outer_grant_valid;
  wire [2:0] trackerList_0_io_outer_grant_bits_addr_beat;
  wire [1:0] trackerList_0_io_outer_grant_bits_client_xact_id;
  wire  trackerList_0_io_outer_grant_bits_manager_xact_id;
  wire  trackerList_0_io_outer_grant_bits_is_builtin_type;
  wire [3:0] trackerList_0_io_outer_grant_bits_g_type;
  wire [63:0] trackerList_0_io_outer_grant_bits_data;
  wire  trackerList_0_io_outer_grant_bits_manager_id;
  wire  trackerList_0_io_outer_finish_ready;
  wire  trackerList_0_io_outer_finish_valid;
  wire  trackerList_0_io_outer_finish_bits_manager_xact_id;
  wire  trackerList_0_io_outer_finish_bits_manager_id;
  wire  trackerList_0_io_alloc_iacq_matches;
  wire  trackerList_0_io_alloc_iacq_can;
  wire  trackerList_0_io_alloc_iacq_should;
  wire  trackerList_0_io_alloc_irel_matches;
  wire  trackerList_0_io_alloc_irel_can;
  wire  trackerList_0_io_alloc_irel_should;
  wire  trackerList_0_io_alloc_oprb_matches;
  wire  trackerList_0_io_alloc_oprb_can;
  wire  trackerList_0_io_alloc_oprb_should;
  wire  trackerList_0_io_alloc_idle;
  wire [25:0] trackerList_0_io_alloc_addr_block;
  wire  trackerList_1_clk;
  wire  trackerList_1_reset;
  wire  trackerList_1_io_inner_acquire_ready;
  wire  trackerList_1_io_inner_acquire_valid;
  wire [25:0] trackerList_1_io_inner_acquire_bits_addr_block;
  wire  trackerList_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] trackerList_1_io_inner_acquire_bits_addr_beat;
  wire  trackerList_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_1_io_inner_acquire_bits_a_type;
  wire [10:0] trackerList_1_io_inner_acquire_bits_union;
  wire [63:0] trackerList_1_io_inner_acquire_bits_data;
  wire  trackerList_1_io_inner_acquire_bits_client_id;
  wire  trackerList_1_io_inner_grant_ready;
  wire  trackerList_1_io_inner_grant_valid;
  wire [2:0] trackerList_1_io_inner_grant_bits_addr_beat;
  wire  trackerList_1_io_inner_grant_bits_client_xact_id;
  wire [1:0] trackerList_1_io_inner_grant_bits_manager_xact_id;
  wire  trackerList_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] trackerList_1_io_inner_grant_bits_g_type;
  wire [63:0] trackerList_1_io_inner_grant_bits_data;
  wire  trackerList_1_io_inner_grant_bits_client_id;
  wire  trackerList_1_io_inner_finish_ready;
  wire  trackerList_1_io_inner_finish_valid;
  wire [1:0] trackerList_1_io_inner_finish_bits_manager_xact_id;
  wire  trackerList_1_io_inner_probe_ready;
  wire  trackerList_1_io_inner_probe_valid;
  wire [25:0] trackerList_1_io_inner_probe_bits_addr_block;
  wire [1:0] trackerList_1_io_inner_probe_bits_p_type;
  wire  trackerList_1_io_inner_probe_bits_client_id;
  wire  trackerList_1_io_inner_release_ready;
  wire  trackerList_1_io_inner_release_valid;
  wire [2:0] trackerList_1_io_inner_release_bits_addr_beat;
  wire [25:0] trackerList_1_io_inner_release_bits_addr_block;
  wire  trackerList_1_io_inner_release_bits_client_xact_id;
  wire  trackerList_1_io_inner_release_bits_voluntary;
  wire [2:0] trackerList_1_io_inner_release_bits_r_type;
  wire [63:0] trackerList_1_io_inner_release_bits_data;
  wire  trackerList_1_io_inner_release_bits_client_id;
  wire  trackerList_1_io_incoherent_0;
  wire  trackerList_1_io_outer_acquire_ready;
  wire  trackerList_1_io_outer_acquire_valid;
  wire [25:0] trackerList_1_io_outer_acquire_bits_addr_block;
  wire [1:0] trackerList_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] trackerList_1_io_outer_acquire_bits_addr_beat;
  wire  trackerList_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_1_io_outer_acquire_bits_a_type;
  wire [10:0] trackerList_1_io_outer_acquire_bits_union;
  wire [63:0] trackerList_1_io_outer_acquire_bits_data;
  wire  trackerList_1_io_outer_probe_ready;
  wire  trackerList_1_io_outer_probe_valid;
  wire [25:0] trackerList_1_io_outer_probe_bits_addr_block;
  wire [1:0] trackerList_1_io_outer_probe_bits_p_type;
  wire  trackerList_1_io_outer_release_ready;
  wire  trackerList_1_io_outer_release_valid;
  wire [2:0] trackerList_1_io_outer_release_bits_addr_beat;
  wire [25:0] trackerList_1_io_outer_release_bits_addr_block;
  wire [1:0] trackerList_1_io_outer_release_bits_client_xact_id;
  wire  trackerList_1_io_outer_release_bits_voluntary;
  wire [2:0] trackerList_1_io_outer_release_bits_r_type;
  wire [63:0] trackerList_1_io_outer_release_bits_data;
  wire  trackerList_1_io_outer_grant_ready;
  wire  trackerList_1_io_outer_grant_valid;
  wire [2:0] trackerList_1_io_outer_grant_bits_addr_beat;
  wire [1:0] trackerList_1_io_outer_grant_bits_client_xact_id;
  wire  trackerList_1_io_outer_grant_bits_manager_xact_id;
  wire  trackerList_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] trackerList_1_io_outer_grant_bits_g_type;
  wire [63:0] trackerList_1_io_outer_grant_bits_data;
  wire  trackerList_1_io_outer_grant_bits_manager_id;
  wire  trackerList_1_io_outer_finish_ready;
  wire  trackerList_1_io_outer_finish_valid;
  wire  trackerList_1_io_outer_finish_bits_manager_xact_id;
  wire  trackerList_1_io_outer_finish_bits_manager_id;
  wire  trackerList_1_io_alloc_iacq_matches;
  wire  trackerList_1_io_alloc_iacq_can;
  wire  trackerList_1_io_alloc_iacq_should;
  wire  trackerList_1_io_alloc_irel_matches;
  wire  trackerList_1_io_alloc_irel_can;
  wire  trackerList_1_io_alloc_irel_should;
  wire  trackerList_1_io_alloc_oprb_matches;
  wire  trackerList_1_io_alloc_oprb_can;
  wire  trackerList_1_io_alloc_oprb_should;
  wire  trackerList_1_io_alloc_idle;
  wire [25:0] trackerList_1_io_alloc_addr_block;
  wire  trackerList_2_clk;
  wire  trackerList_2_reset;
  wire  trackerList_2_io_inner_acquire_ready;
  wire  trackerList_2_io_inner_acquire_valid;
  wire [25:0] trackerList_2_io_inner_acquire_bits_addr_block;
  wire  trackerList_2_io_inner_acquire_bits_client_xact_id;
  wire [2:0] trackerList_2_io_inner_acquire_bits_addr_beat;
  wire  trackerList_2_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_2_io_inner_acquire_bits_a_type;
  wire [10:0] trackerList_2_io_inner_acquire_bits_union;
  wire [63:0] trackerList_2_io_inner_acquire_bits_data;
  wire  trackerList_2_io_inner_acquire_bits_client_id;
  wire  trackerList_2_io_inner_grant_ready;
  wire  trackerList_2_io_inner_grant_valid;
  wire [2:0] trackerList_2_io_inner_grant_bits_addr_beat;
  wire  trackerList_2_io_inner_grant_bits_client_xact_id;
  wire [1:0] trackerList_2_io_inner_grant_bits_manager_xact_id;
  wire  trackerList_2_io_inner_grant_bits_is_builtin_type;
  wire [3:0] trackerList_2_io_inner_grant_bits_g_type;
  wire [63:0] trackerList_2_io_inner_grant_bits_data;
  wire  trackerList_2_io_inner_grant_bits_client_id;
  wire  trackerList_2_io_inner_finish_ready;
  wire  trackerList_2_io_inner_finish_valid;
  wire [1:0] trackerList_2_io_inner_finish_bits_manager_xact_id;
  wire  trackerList_2_io_inner_probe_ready;
  wire  trackerList_2_io_inner_probe_valid;
  wire [25:0] trackerList_2_io_inner_probe_bits_addr_block;
  wire [1:0] trackerList_2_io_inner_probe_bits_p_type;
  wire  trackerList_2_io_inner_probe_bits_client_id;
  wire  trackerList_2_io_inner_release_ready;
  wire  trackerList_2_io_inner_release_valid;
  wire [2:0] trackerList_2_io_inner_release_bits_addr_beat;
  wire [25:0] trackerList_2_io_inner_release_bits_addr_block;
  wire  trackerList_2_io_inner_release_bits_client_xact_id;
  wire  trackerList_2_io_inner_release_bits_voluntary;
  wire [2:0] trackerList_2_io_inner_release_bits_r_type;
  wire [63:0] trackerList_2_io_inner_release_bits_data;
  wire  trackerList_2_io_inner_release_bits_client_id;
  wire  trackerList_2_io_incoherent_0;
  wire  trackerList_2_io_outer_acquire_ready;
  wire  trackerList_2_io_outer_acquire_valid;
  wire [25:0] trackerList_2_io_outer_acquire_bits_addr_block;
  wire [1:0] trackerList_2_io_outer_acquire_bits_client_xact_id;
  wire [2:0] trackerList_2_io_outer_acquire_bits_addr_beat;
  wire  trackerList_2_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_2_io_outer_acquire_bits_a_type;
  wire [10:0] trackerList_2_io_outer_acquire_bits_union;
  wire [63:0] trackerList_2_io_outer_acquire_bits_data;
  wire  trackerList_2_io_outer_probe_ready;
  wire  trackerList_2_io_outer_probe_valid;
  wire [25:0] trackerList_2_io_outer_probe_bits_addr_block;
  wire [1:0] trackerList_2_io_outer_probe_bits_p_type;
  wire  trackerList_2_io_outer_release_ready;
  wire  trackerList_2_io_outer_release_valid;
  wire [2:0] trackerList_2_io_outer_release_bits_addr_beat;
  wire [25:0] trackerList_2_io_outer_release_bits_addr_block;
  wire [1:0] trackerList_2_io_outer_release_bits_client_xact_id;
  wire  trackerList_2_io_outer_release_bits_voluntary;
  wire [2:0] trackerList_2_io_outer_release_bits_r_type;
  wire [63:0] trackerList_2_io_outer_release_bits_data;
  wire  trackerList_2_io_outer_grant_ready;
  wire  trackerList_2_io_outer_grant_valid;
  wire [2:0] trackerList_2_io_outer_grant_bits_addr_beat;
  wire [1:0] trackerList_2_io_outer_grant_bits_client_xact_id;
  wire  trackerList_2_io_outer_grant_bits_manager_xact_id;
  wire  trackerList_2_io_outer_grant_bits_is_builtin_type;
  wire [3:0] trackerList_2_io_outer_grant_bits_g_type;
  wire [63:0] trackerList_2_io_outer_grant_bits_data;
  wire  trackerList_2_io_outer_grant_bits_manager_id;
  wire  trackerList_2_io_outer_finish_ready;
  wire  trackerList_2_io_outer_finish_valid;
  wire  trackerList_2_io_outer_finish_bits_manager_xact_id;
  wire  trackerList_2_io_outer_finish_bits_manager_id;
  wire  trackerList_2_io_alloc_iacq_matches;
  wire  trackerList_2_io_alloc_iacq_can;
  wire  trackerList_2_io_alloc_iacq_should;
  wire  trackerList_2_io_alloc_irel_matches;
  wire  trackerList_2_io_alloc_irel_can;
  wire  trackerList_2_io_alloc_irel_should;
  wire  trackerList_2_io_alloc_oprb_matches;
  wire  trackerList_2_io_alloc_oprb_can;
  wire  trackerList_2_io_alloc_oprb_should;
  wire  trackerList_2_io_alloc_idle;
  wire [25:0] trackerList_2_io_alloc_addr_block;
  wire  outer_arb_clk;
  wire  outer_arb_reset;
  wire  outer_arb_io_in_0_acquire_ready;
  wire  outer_arb_io_in_0_acquire_valid;
  wire [25:0] outer_arb_io_in_0_acquire_bits_addr_block;
  wire [1:0] outer_arb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_0_acquire_bits_addr_beat;
  wire  outer_arb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_0_acquire_bits_a_type;
  wire [10:0] outer_arb_io_in_0_acquire_bits_union;
  wire [63:0] outer_arb_io_in_0_acquire_bits_data;
  wire  outer_arb_io_in_0_probe_ready;
  wire  outer_arb_io_in_0_probe_valid;
  wire [25:0] outer_arb_io_in_0_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_0_probe_bits_p_type;
  wire  outer_arb_io_in_0_release_ready;
  wire  outer_arb_io_in_0_release_valid;
  wire [2:0] outer_arb_io_in_0_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_0_release_bits_addr_block;
  wire [1:0] outer_arb_io_in_0_release_bits_client_xact_id;
  wire  outer_arb_io_in_0_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_0_release_bits_r_type;
  wire [63:0] outer_arb_io_in_0_release_bits_data;
  wire  outer_arb_io_in_0_grant_ready;
  wire  outer_arb_io_in_0_grant_valid;
  wire [2:0] outer_arb_io_in_0_grant_bits_addr_beat;
  wire [1:0] outer_arb_io_in_0_grant_bits_client_xact_id;
  wire  outer_arb_io_in_0_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_0_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_0_grant_bits_data;
  wire  outer_arb_io_in_0_grant_bits_manager_id;
  wire  outer_arb_io_in_0_finish_ready;
  wire  outer_arb_io_in_0_finish_valid;
  wire  outer_arb_io_in_0_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_0_finish_bits_manager_id;
  wire  outer_arb_io_in_1_acquire_ready;
  wire  outer_arb_io_in_1_acquire_valid;
  wire [25:0] outer_arb_io_in_1_acquire_bits_addr_block;
  wire [1:0] outer_arb_io_in_1_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_1_acquire_bits_addr_beat;
  wire  outer_arb_io_in_1_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_1_acquire_bits_a_type;
  wire [10:0] outer_arb_io_in_1_acquire_bits_union;
  wire [63:0] outer_arb_io_in_1_acquire_bits_data;
  wire  outer_arb_io_in_1_probe_ready;
  wire  outer_arb_io_in_1_probe_valid;
  wire [25:0] outer_arb_io_in_1_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_1_probe_bits_p_type;
  wire  outer_arb_io_in_1_release_ready;
  wire  outer_arb_io_in_1_release_valid;
  wire [2:0] outer_arb_io_in_1_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_1_release_bits_addr_block;
  wire [1:0] outer_arb_io_in_1_release_bits_client_xact_id;
  wire  outer_arb_io_in_1_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_1_release_bits_r_type;
  wire [63:0] outer_arb_io_in_1_release_bits_data;
  wire  outer_arb_io_in_1_grant_ready;
  wire  outer_arb_io_in_1_grant_valid;
  wire [2:0] outer_arb_io_in_1_grant_bits_addr_beat;
  wire [1:0] outer_arb_io_in_1_grant_bits_client_xact_id;
  wire  outer_arb_io_in_1_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_1_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_1_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_1_grant_bits_data;
  wire  outer_arb_io_in_1_grant_bits_manager_id;
  wire  outer_arb_io_in_1_finish_ready;
  wire  outer_arb_io_in_1_finish_valid;
  wire  outer_arb_io_in_1_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_1_finish_bits_manager_id;
  wire  outer_arb_io_in_2_acquire_ready;
  wire  outer_arb_io_in_2_acquire_valid;
  wire [25:0] outer_arb_io_in_2_acquire_bits_addr_block;
  wire [1:0] outer_arb_io_in_2_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_2_acquire_bits_addr_beat;
  wire  outer_arb_io_in_2_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_2_acquire_bits_a_type;
  wire [10:0] outer_arb_io_in_2_acquire_bits_union;
  wire [63:0] outer_arb_io_in_2_acquire_bits_data;
  wire  outer_arb_io_in_2_probe_ready;
  wire  outer_arb_io_in_2_probe_valid;
  wire [25:0] outer_arb_io_in_2_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_2_probe_bits_p_type;
  wire  outer_arb_io_in_2_release_ready;
  wire  outer_arb_io_in_2_release_valid;
  wire [2:0] outer_arb_io_in_2_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_2_release_bits_addr_block;
  wire [1:0] outer_arb_io_in_2_release_bits_client_xact_id;
  wire  outer_arb_io_in_2_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_2_release_bits_r_type;
  wire [63:0] outer_arb_io_in_2_release_bits_data;
  wire  outer_arb_io_in_2_grant_ready;
  wire  outer_arb_io_in_2_grant_valid;
  wire [2:0] outer_arb_io_in_2_grant_bits_addr_beat;
  wire [1:0] outer_arb_io_in_2_grant_bits_client_xact_id;
  wire  outer_arb_io_in_2_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_2_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_2_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_2_grant_bits_data;
  wire  outer_arb_io_in_2_grant_bits_manager_id;
  wire  outer_arb_io_in_2_finish_ready;
  wire  outer_arb_io_in_2_finish_valid;
  wire  outer_arb_io_in_2_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_2_finish_bits_manager_id;
  wire  outer_arb_io_out_acquire_ready;
  wire  outer_arb_io_out_acquire_valid;
  wire [25:0] outer_arb_io_out_acquire_bits_addr_block;
  wire [1:0] outer_arb_io_out_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_out_acquire_bits_addr_beat;
  wire  outer_arb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_out_acquire_bits_a_type;
  wire [10:0] outer_arb_io_out_acquire_bits_union;
  wire [63:0] outer_arb_io_out_acquire_bits_data;
  wire  outer_arb_io_out_probe_ready;
  wire  outer_arb_io_out_probe_valid;
  wire [25:0] outer_arb_io_out_probe_bits_addr_block;
  wire [1:0] outer_arb_io_out_probe_bits_p_type;
  wire  outer_arb_io_out_release_ready;
  wire  outer_arb_io_out_release_valid;
  wire [2:0] outer_arb_io_out_release_bits_addr_beat;
  wire [25:0] outer_arb_io_out_release_bits_addr_block;
  wire [1:0] outer_arb_io_out_release_bits_client_xact_id;
  wire  outer_arb_io_out_release_bits_voluntary;
  wire [2:0] outer_arb_io_out_release_bits_r_type;
  wire [63:0] outer_arb_io_out_release_bits_data;
  wire  outer_arb_io_out_grant_ready;
  wire  outer_arb_io_out_grant_valid;
  wire [2:0] outer_arb_io_out_grant_bits_addr_beat;
  wire [1:0] outer_arb_io_out_grant_bits_client_xact_id;
  wire  outer_arb_io_out_grant_bits_manager_xact_id;
  wire  outer_arb_io_out_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_out_grant_bits_g_type;
  wire [63:0] outer_arb_io_out_grant_bits_data;
  wire  outer_arb_io_out_grant_bits_manager_id;
  wire  outer_arb_io_out_finish_ready;
  wire  outer_arb_io_out_finish_valid;
  wire  outer_arb_io_out_finish_bits_manager_xact_id;
  wire  outer_arb_io_out_finish_bits_manager_id;
  wire  T_1215;
  wire  T_1216;
  wire  irel_vs_iacq_conflict;
  wire  T_1218;
  wire [1:0] T_1219;
  wire [2:0] T_1220;
  wire [1:0] T_1221;
  wire [2:0] T_1222;
  wire  T_1223;
  wire  T_1224;
  wire  T_1225;
  wire [2:0] T_1231;
  wire [2:0] T_1232;
  wire [2:0] T_1233;
  wire [1:0] T_1234;
  wire [2:0] T_1235;
  wire  T_1237;
  wire  T_1239;
  wire [2:0] T_1241;
  wire [2:0] T_1242;
  wire  T_1244;
  wire  T_1245;
  wire  T_1248;
  wire  T_1249;
  wire  T_1250;
  wire  T_1251;
  wire  T_1254;
  wire  T_1255;
  wire  T_1256;
  wire  T_1259;
  wire  T_1260;
  wire  T_1261;
  wire [1:0] T_1262;
  wire [2:0] T_1263;
  wire [1:0] T_1264;
  wire [2:0] T_1265;
  wire  T_1266;
  wire  T_1267;
  wire  T_1268;
  wire [2:0] T_1274;
  wire [2:0] T_1275;
  wire [2:0] T_1276;
  wire [1:0] T_1277;
  wire [2:0] T_1278;
  wire  T_1280;
  wire  T_1282;
  wire [2:0] T_1285;
  wire [2:0] T_1286;
  wire  T_1288;
  wire  T_1293;
  wire  T_1294;
  wire  T_1298;
  wire  T_1299;
  wire  T_1303;
  wire  T_1304;
  wire  LockingRRArbiter_7_1_clk;
  wire  LockingRRArbiter_7_1_reset;
  wire  LockingRRArbiter_7_1_io_in_0_ready;
  wire  LockingRRArbiter_7_1_io_in_0_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_0_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_0_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_0_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_1_ready;
  wire  LockingRRArbiter_7_1_io_in_1_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_1_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_1_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_1_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_2_ready;
  wire  LockingRRArbiter_7_1_io_in_2_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_2_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_2_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_2_bits_client_id;
  wire  LockingRRArbiter_7_1_io_out_ready;
  wire  LockingRRArbiter_7_1_io_out_valid;
  wire [25:0] LockingRRArbiter_7_1_io_out_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_out_bits_p_type;
  wire  LockingRRArbiter_7_1_io_out_bits_client_id;
  wire [1:0] LockingRRArbiter_7_1_io_chosen;
  wire  LockingRRArbiter_8_1_clk;
  wire  LockingRRArbiter_8_1_reset;
  wire  LockingRRArbiter_8_1_io_in_0_ready;
  wire  LockingRRArbiter_8_1_io_in_0_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_0_bits_addr_beat;
  wire  LockingRRArbiter_8_1_io_in_0_bits_client_xact_id;
  wire [1:0] LockingRRArbiter_8_1_io_in_0_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_0_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_0_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_0_bits_data;
  wire  LockingRRArbiter_8_1_io_in_0_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_1_ready;
  wire  LockingRRArbiter_8_1_io_in_1_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_1_bits_addr_beat;
  wire  LockingRRArbiter_8_1_io_in_1_bits_client_xact_id;
  wire [1:0] LockingRRArbiter_8_1_io_in_1_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_1_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_1_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_1_bits_data;
  wire  LockingRRArbiter_8_1_io_in_1_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_2_ready;
  wire  LockingRRArbiter_8_1_io_in_2_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_2_bits_addr_beat;
  wire  LockingRRArbiter_8_1_io_in_2_bits_client_xact_id;
  wire [1:0] LockingRRArbiter_8_1_io_in_2_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_2_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_2_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_2_bits_data;
  wire  LockingRRArbiter_8_1_io_in_2_bits_client_id;
  wire  LockingRRArbiter_8_1_io_out_ready;
  wire  LockingRRArbiter_8_1_io_out_valid;
  wire [2:0] LockingRRArbiter_8_1_io_out_bits_addr_beat;
  wire  LockingRRArbiter_8_1_io_out_bits_client_xact_id;
  wire [1:0] LockingRRArbiter_8_1_io_out_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_out_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_out_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_out_bits_data;
  wire  LockingRRArbiter_8_1_io_out_bits_client_id;
  wire [1:0] LockingRRArbiter_8_1_io_chosen;
  wire  T_1307;
  wire  T_1308;
  wire  T_1310;
  wire  T_1311;
  wire  T_1313;
  wire  T_1314;
  wire [1:0] T_1316;
  wire  T_1318;
  wire  T_1322;
  wire  T_1323;
  wire  T_1324;
  wire  T_1328;
  wire  T_1329;
  wire  T_1331;
  wire  GEN_0;
  reg [31:0] GEN_3;
  wire  GEN_1;
  reg [31:0] GEN_4;
  wire  GEN_2;
  reg [31:0] GEN_5;
  BufferedBroadcastVoluntaryReleaseTracker trackerList_0 (
    .clk(trackerList_0_clk),
    .reset(trackerList_0_reset),
    .io_inner_acquire_ready(trackerList_0_io_inner_acquire_ready),
    .io_inner_acquire_valid(trackerList_0_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(trackerList_0_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(trackerList_0_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(trackerList_0_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(trackerList_0_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(trackerList_0_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(trackerList_0_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(trackerList_0_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(trackerList_0_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(trackerList_0_io_inner_grant_ready),
    .io_inner_grant_valid(trackerList_0_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(trackerList_0_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(trackerList_0_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(trackerList_0_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(trackerList_0_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(trackerList_0_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(trackerList_0_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(trackerList_0_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(trackerList_0_io_inner_finish_ready),
    .io_inner_finish_valid(trackerList_0_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(trackerList_0_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(trackerList_0_io_inner_probe_ready),
    .io_inner_probe_valid(trackerList_0_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(trackerList_0_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(trackerList_0_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(trackerList_0_io_inner_probe_bits_client_id),
    .io_inner_release_ready(trackerList_0_io_inner_release_ready),
    .io_inner_release_valid(trackerList_0_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(trackerList_0_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(trackerList_0_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(trackerList_0_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(trackerList_0_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(trackerList_0_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(trackerList_0_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(trackerList_0_io_inner_release_bits_client_id),
    .io_incoherent_0(trackerList_0_io_incoherent_0),
    .io_outer_acquire_ready(trackerList_0_io_outer_acquire_ready),
    .io_outer_acquire_valid(trackerList_0_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(trackerList_0_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(trackerList_0_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(trackerList_0_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(trackerList_0_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(trackerList_0_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(trackerList_0_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(trackerList_0_io_outer_acquire_bits_data),
    .io_outer_probe_ready(trackerList_0_io_outer_probe_ready),
    .io_outer_probe_valid(trackerList_0_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(trackerList_0_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(trackerList_0_io_outer_probe_bits_p_type),
    .io_outer_release_ready(trackerList_0_io_outer_release_ready),
    .io_outer_release_valid(trackerList_0_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(trackerList_0_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(trackerList_0_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(trackerList_0_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(trackerList_0_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(trackerList_0_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(trackerList_0_io_outer_release_bits_data),
    .io_outer_grant_ready(trackerList_0_io_outer_grant_ready),
    .io_outer_grant_valid(trackerList_0_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(trackerList_0_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(trackerList_0_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(trackerList_0_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(trackerList_0_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(trackerList_0_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(trackerList_0_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(trackerList_0_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(trackerList_0_io_outer_finish_ready),
    .io_outer_finish_valid(trackerList_0_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(trackerList_0_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(trackerList_0_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(trackerList_0_io_alloc_iacq_matches),
    .io_alloc_iacq_can(trackerList_0_io_alloc_iacq_can),
    .io_alloc_iacq_should(trackerList_0_io_alloc_iacq_should),
    .io_alloc_irel_matches(trackerList_0_io_alloc_irel_matches),
    .io_alloc_irel_can(trackerList_0_io_alloc_irel_can),
    .io_alloc_irel_should(trackerList_0_io_alloc_irel_should),
    .io_alloc_oprb_matches(trackerList_0_io_alloc_oprb_matches),
    .io_alloc_oprb_can(trackerList_0_io_alloc_oprb_can),
    .io_alloc_oprb_should(trackerList_0_io_alloc_oprb_should),
    .io_alloc_idle(trackerList_0_io_alloc_idle),
    .io_alloc_addr_block(trackerList_0_io_alloc_addr_block)
  );
  BufferedBroadcastAcquireTracker trackerList_1 (
    .clk(trackerList_1_clk),
    .reset(trackerList_1_reset),
    .io_inner_acquire_ready(trackerList_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(trackerList_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(trackerList_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(trackerList_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(trackerList_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(trackerList_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(trackerList_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(trackerList_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(trackerList_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(trackerList_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(trackerList_1_io_inner_grant_ready),
    .io_inner_grant_valid(trackerList_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(trackerList_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(trackerList_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(trackerList_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(trackerList_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(trackerList_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(trackerList_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(trackerList_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(trackerList_1_io_inner_finish_ready),
    .io_inner_finish_valid(trackerList_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(trackerList_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(trackerList_1_io_inner_probe_ready),
    .io_inner_probe_valid(trackerList_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(trackerList_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(trackerList_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(trackerList_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(trackerList_1_io_inner_release_ready),
    .io_inner_release_valid(trackerList_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(trackerList_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(trackerList_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(trackerList_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(trackerList_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(trackerList_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(trackerList_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(trackerList_1_io_inner_release_bits_client_id),
    .io_incoherent_0(trackerList_1_io_incoherent_0),
    .io_outer_acquire_ready(trackerList_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(trackerList_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(trackerList_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(trackerList_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(trackerList_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(trackerList_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(trackerList_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(trackerList_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(trackerList_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(trackerList_1_io_outer_probe_ready),
    .io_outer_probe_valid(trackerList_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(trackerList_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(trackerList_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(trackerList_1_io_outer_release_ready),
    .io_outer_release_valid(trackerList_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(trackerList_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(trackerList_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(trackerList_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(trackerList_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(trackerList_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(trackerList_1_io_outer_release_bits_data),
    .io_outer_grant_ready(trackerList_1_io_outer_grant_ready),
    .io_outer_grant_valid(trackerList_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(trackerList_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(trackerList_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(trackerList_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(trackerList_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(trackerList_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(trackerList_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(trackerList_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(trackerList_1_io_outer_finish_ready),
    .io_outer_finish_valid(trackerList_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(trackerList_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(trackerList_1_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(trackerList_1_io_alloc_iacq_matches),
    .io_alloc_iacq_can(trackerList_1_io_alloc_iacq_can),
    .io_alloc_iacq_should(trackerList_1_io_alloc_iacq_should),
    .io_alloc_irel_matches(trackerList_1_io_alloc_irel_matches),
    .io_alloc_irel_can(trackerList_1_io_alloc_irel_can),
    .io_alloc_irel_should(trackerList_1_io_alloc_irel_should),
    .io_alloc_oprb_matches(trackerList_1_io_alloc_oprb_matches),
    .io_alloc_oprb_can(trackerList_1_io_alloc_oprb_can),
    .io_alloc_oprb_should(trackerList_1_io_alloc_oprb_should),
    .io_alloc_idle(trackerList_1_io_alloc_idle),
    .io_alloc_addr_block(trackerList_1_io_alloc_addr_block)
  );
  BufferedBroadcastAcquireTracker_1 trackerList_2 (
    .clk(trackerList_2_clk),
    .reset(trackerList_2_reset),
    .io_inner_acquire_ready(trackerList_2_io_inner_acquire_ready),
    .io_inner_acquire_valid(trackerList_2_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(trackerList_2_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(trackerList_2_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(trackerList_2_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(trackerList_2_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(trackerList_2_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(trackerList_2_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(trackerList_2_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(trackerList_2_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(trackerList_2_io_inner_grant_ready),
    .io_inner_grant_valid(trackerList_2_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(trackerList_2_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(trackerList_2_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(trackerList_2_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(trackerList_2_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(trackerList_2_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(trackerList_2_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(trackerList_2_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(trackerList_2_io_inner_finish_ready),
    .io_inner_finish_valid(trackerList_2_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(trackerList_2_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(trackerList_2_io_inner_probe_ready),
    .io_inner_probe_valid(trackerList_2_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(trackerList_2_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(trackerList_2_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(trackerList_2_io_inner_probe_bits_client_id),
    .io_inner_release_ready(trackerList_2_io_inner_release_ready),
    .io_inner_release_valid(trackerList_2_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(trackerList_2_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(trackerList_2_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(trackerList_2_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(trackerList_2_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(trackerList_2_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(trackerList_2_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(trackerList_2_io_inner_release_bits_client_id),
    .io_incoherent_0(trackerList_2_io_incoherent_0),
    .io_outer_acquire_ready(trackerList_2_io_outer_acquire_ready),
    .io_outer_acquire_valid(trackerList_2_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(trackerList_2_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(trackerList_2_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(trackerList_2_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(trackerList_2_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(trackerList_2_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(trackerList_2_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(trackerList_2_io_outer_acquire_bits_data),
    .io_outer_probe_ready(trackerList_2_io_outer_probe_ready),
    .io_outer_probe_valid(trackerList_2_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(trackerList_2_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(trackerList_2_io_outer_probe_bits_p_type),
    .io_outer_release_ready(trackerList_2_io_outer_release_ready),
    .io_outer_release_valid(trackerList_2_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(trackerList_2_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(trackerList_2_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(trackerList_2_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(trackerList_2_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(trackerList_2_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(trackerList_2_io_outer_release_bits_data),
    .io_outer_grant_ready(trackerList_2_io_outer_grant_ready),
    .io_outer_grant_valid(trackerList_2_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(trackerList_2_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(trackerList_2_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(trackerList_2_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(trackerList_2_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(trackerList_2_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(trackerList_2_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(trackerList_2_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(trackerList_2_io_outer_finish_ready),
    .io_outer_finish_valid(trackerList_2_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(trackerList_2_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(trackerList_2_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(trackerList_2_io_alloc_iacq_matches),
    .io_alloc_iacq_can(trackerList_2_io_alloc_iacq_can),
    .io_alloc_iacq_should(trackerList_2_io_alloc_iacq_should),
    .io_alloc_irel_matches(trackerList_2_io_alloc_irel_matches),
    .io_alloc_irel_can(trackerList_2_io_alloc_irel_can),
    .io_alloc_irel_should(trackerList_2_io_alloc_irel_should),
    .io_alloc_oprb_matches(trackerList_2_io_alloc_oprb_matches),
    .io_alloc_oprb_can(trackerList_2_io_alloc_oprb_can),
    .io_alloc_oprb_should(trackerList_2_io_alloc_oprb_should),
    .io_alloc_idle(trackerList_2_io_alloc_idle),
    .io_alloc_addr_block(trackerList_2_io_alloc_addr_block)
  );
  ClientTileLinkIOArbiter outer_arb (
    .clk(outer_arb_clk),
    .reset(outer_arb_reset),
    .io_in_0_acquire_ready(outer_arb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(outer_arb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(outer_arb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(outer_arb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(outer_arb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(outer_arb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(outer_arb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(outer_arb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(outer_arb_io_in_0_acquire_bits_data),
    .io_in_0_probe_ready(outer_arb_io_in_0_probe_ready),
    .io_in_0_probe_valid(outer_arb_io_in_0_probe_valid),
    .io_in_0_probe_bits_addr_block(outer_arb_io_in_0_probe_bits_addr_block),
    .io_in_0_probe_bits_p_type(outer_arb_io_in_0_probe_bits_p_type),
    .io_in_0_release_ready(outer_arb_io_in_0_release_ready),
    .io_in_0_release_valid(outer_arb_io_in_0_release_valid),
    .io_in_0_release_bits_addr_beat(outer_arb_io_in_0_release_bits_addr_beat),
    .io_in_0_release_bits_addr_block(outer_arb_io_in_0_release_bits_addr_block),
    .io_in_0_release_bits_client_xact_id(outer_arb_io_in_0_release_bits_client_xact_id),
    .io_in_0_release_bits_voluntary(outer_arb_io_in_0_release_bits_voluntary),
    .io_in_0_release_bits_r_type(outer_arb_io_in_0_release_bits_r_type),
    .io_in_0_release_bits_data(outer_arb_io_in_0_release_bits_data),
    .io_in_0_grant_ready(outer_arb_io_in_0_grant_ready),
    .io_in_0_grant_valid(outer_arb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(outer_arb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(outer_arb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(outer_arb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(outer_arb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(outer_arb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(outer_arb_io_in_0_grant_bits_data),
    .io_in_0_grant_bits_manager_id(outer_arb_io_in_0_grant_bits_manager_id),
    .io_in_0_finish_ready(outer_arb_io_in_0_finish_ready),
    .io_in_0_finish_valid(outer_arb_io_in_0_finish_valid),
    .io_in_0_finish_bits_manager_xact_id(outer_arb_io_in_0_finish_bits_manager_xact_id),
    .io_in_0_finish_bits_manager_id(outer_arb_io_in_0_finish_bits_manager_id),
    .io_in_1_acquire_ready(outer_arb_io_in_1_acquire_ready),
    .io_in_1_acquire_valid(outer_arb_io_in_1_acquire_valid),
    .io_in_1_acquire_bits_addr_block(outer_arb_io_in_1_acquire_bits_addr_block),
    .io_in_1_acquire_bits_client_xact_id(outer_arb_io_in_1_acquire_bits_client_xact_id),
    .io_in_1_acquire_bits_addr_beat(outer_arb_io_in_1_acquire_bits_addr_beat),
    .io_in_1_acquire_bits_is_builtin_type(outer_arb_io_in_1_acquire_bits_is_builtin_type),
    .io_in_1_acquire_bits_a_type(outer_arb_io_in_1_acquire_bits_a_type),
    .io_in_1_acquire_bits_union(outer_arb_io_in_1_acquire_bits_union),
    .io_in_1_acquire_bits_data(outer_arb_io_in_1_acquire_bits_data),
    .io_in_1_probe_ready(outer_arb_io_in_1_probe_ready),
    .io_in_1_probe_valid(outer_arb_io_in_1_probe_valid),
    .io_in_1_probe_bits_addr_block(outer_arb_io_in_1_probe_bits_addr_block),
    .io_in_1_probe_bits_p_type(outer_arb_io_in_1_probe_bits_p_type),
    .io_in_1_release_ready(outer_arb_io_in_1_release_ready),
    .io_in_1_release_valid(outer_arb_io_in_1_release_valid),
    .io_in_1_release_bits_addr_beat(outer_arb_io_in_1_release_bits_addr_beat),
    .io_in_1_release_bits_addr_block(outer_arb_io_in_1_release_bits_addr_block),
    .io_in_1_release_bits_client_xact_id(outer_arb_io_in_1_release_bits_client_xact_id),
    .io_in_1_release_bits_voluntary(outer_arb_io_in_1_release_bits_voluntary),
    .io_in_1_release_bits_r_type(outer_arb_io_in_1_release_bits_r_type),
    .io_in_1_release_bits_data(outer_arb_io_in_1_release_bits_data),
    .io_in_1_grant_ready(outer_arb_io_in_1_grant_ready),
    .io_in_1_grant_valid(outer_arb_io_in_1_grant_valid),
    .io_in_1_grant_bits_addr_beat(outer_arb_io_in_1_grant_bits_addr_beat),
    .io_in_1_grant_bits_client_xact_id(outer_arb_io_in_1_grant_bits_client_xact_id),
    .io_in_1_grant_bits_manager_xact_id(outer_arb_io_in_1_grant_bits_manager_xact_id),
    .io_in_1_grant_bits_is_builtin_type(outer_arb_io_in_1_grant_bits_is_builtin_type),
    .io_in_1_grant_bits_g_type(outer_arb_io_in_1_grant_bits_g_type),
    .io_in_1_grant_bits_data(outer_arb_io_in_1_grant_bits_data),
    .io_in_1_grant_bits_manager_id(outer_arb_io_in_1_grant_bits_manager_id),
    .io_in_1_finish_ready(outer_arb_io_in_1_finish_ready),
    .io_in_1_finish_valid(outer_arb_io_in_1_finish_valid),
    .io_in_1_finish_bits_manager_xact_id(outer_arb_io_in_1_finish_bits_manager_xact_id),
    .io_in_1_finish_bits_manager_id(outer_arb_io_in_1_finish_bits_manager_id),
    .io_in_2_acquire_ready(outer_arb_io_in_2_acquire_ready),
    .io_in_2_acquire_valid(outer_arb_io_in_2_acquire_valid),
    .io_in_2_acquire_bits_addr_block(outer_arb_io_in_2_acquire_bits_addr_block),
    .io_in_2_acquire_bits_client_xact_id(outer_arb_io_in_2_acquire_bits_client_xact_id),
    .io_in_2_acquire_bits_addr_beat(outer_arb_io_in_2_acquire_bits_addr_beat),
    .io_in_2_acquire_bits_is_builtin_type(outer_arb_io_in_2_acquire_bits_is_builtin_type),
    .io_in_2_acquire_bits_a_type(outer_arb_io_in_2_acquire_bits_a_type),
    .io_in_2_acquire_bits_union(outer_arb_io_in_2_acquire_bits_union),
    .io_in_2_acquire_bits_data(outer_arb_io_in_2_acquire_bits_data),
    .io_in_2_probe_ready(outer_arb_io_in_2_probe_ready),
    .io_in_2_probe_valid(outer_arb_io_in_2_probe_valid),
    .io_in_2_probe_bits_addr_block(outer_arb_io_in_2_probe_bits_addr_block),
    .io_in_2_probe_bits_p_type(outer_arb_io_in_2_probe_bits_p_type),
    .io_in_2_release_ready(outer_arb_io_in_2_release_ready),
    .io_in_2_release_valid(outer_arb_io_in_2_release_valid),
    .io_in_2_release_bits_addr_beat(outer_arb_io_in_2_release_bits_addr_beat),
    .io_in_2_release_bits_addr_block(outer_arb_io_in_2_release_bits_addr_block),
    .io_in_2_release_bits_client_xact_id(outer_arb_io_in_2_release_bits_client_xact_id),
    .io_in_2_release_bits_voluntary(outer_arb_io_in_2_release_bits_voluntary),
    .io_in_2_release_bits_r_type(outer_arb_io_in_2_release_bits_r_type),
    .io_in_2_release_bits_data(outer_arb_io_in_2_release_bits_data),
    .io_in_2_grant_ready(outer_arb_io_in_2_grant_ready),
    .io_in_2_grant_valid(outer_arb_io_in_2_grant_valid),
    .io_in_2_grant_bits_addr_beat(outer_arb_io_in_2_grant_bits_addr_beat),
    .io_in_2_grant_bits_client_xact_id(outer_arb_io_in_2_grant_bits_client_xact_id),
    .io_in_2_grant_bits_manager_xact_id(outer_arb_io_in_2_grant_bits_manager_xact_id),
    .io_in_2_grant_bits_is_builtin_type(outer_arb_io_in_2_grant_bits_is_builtin_type),
    .io_in_2_grant_bits_g_type(outer_arb_io_in_2_grant_bits_g_type),
    .io_in_2_grant_bits_data(outer_arb_io_in_2_grant_bits_data),
    .io_in_2_grant_bits_manager_id(outer_arb_io_in_2_grant_bits_manager_id),
    .io_in_2_finish_ready(outer_arb_io_in_2_finish_ready),
    .io_in_2_finish_valid(outer_arb_io_in_2_finish_valid),
    .io_in_2_finish_bits_manager_xact_id(outer_arb_io_in_2_finish_bits_manager_xact_id),
    .io_in_2_finish_bits_manager_id(outer_arb_io_in_2_finish_bits_manager_id),
    .io_out_acquire_ready(outer_arb_io_out_acquire_ready),
    .io_out_acquire_valid(outer_arb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(outer_arb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(outer_arb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(outer_arb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(outer_arb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(outer_arb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(outer_arb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(outer_arb_io_out_acquire_bits_data),
    .io_out_probe_ready(outer_arb_io_out_probe_ready),
    .io_out_probe_valid(outer_arb_io_out_probe_valid),
    .io_out_probe_bits_addr_block(outer_arb_io_out_probe_bits_addr_block),
    .io_out_probe_bits_p_type(outer_arb_io_out_probe_bits_p_type),
    .io_out_release_ready(outer_arb_io_out_release_ready),
    .io_out_release_valid(outer_arb_io_out_release_valid),
    .io_out_release_bits_addr_beat(outer_arb_io_out_release_bits_addr_beat),
    .io_out_release_bits_addr_block(outer_arb_io_out_release_bits_addr_block),
    .io_out_release_bits_client_xact_id(outer_arb_io_out_release_bits_client_xact_id),
    .io_out_release_bits_voluntary(outer_arb_io_out_release_bits_voluntary),
    .io_out_release_bits_r_type(outer_arb_io_out_release_bits_r_type),
    .io_out_release_bits_data(outer_arb_io_out_release_bits_data),
    .io_out_grant_ready(outer_arb_io_out_grant_ready),
    .io_out_grant_valid(outer_arb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(outer_arb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(outer_arb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(outer_arb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(outer_arb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(outer_arb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(outer_arb_io_out_grant_bits_data),
    .io_out_grant_bits_manager_id(outer_arb_io_out_grant_bits_manager_id),
    .io_out_finish_ready(outer_arb_io_out_finish_ready),
    .io_out_finish_valid(outer_arb_io_out_finish_valid),
    .io_out_finish_bits_manager_xact_id(outer_arb_io_out_finish_bits_manager_xact_id),
    .io_out_finish_bits_manager_id(outer_arb_io_out_finish_bits_manager_id)
  );
  LockingRRArbiter_7 LockingRRArbiter_7_1 (
    .clk(LockingRRArbiter_7_1_clk),
    .reset(LockingRRArbiter_7_1_reset),
    .io_in_0_ready(LockingRRArbiter_7_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_7_1_io_in_0_valid),
    .io_in_0_bits_addr_block(LockingRRArbiter_7_1_io_in_0_bits_addr_block),
    .io_in_0_bits_p_type(LockingRRArbiter_7_1_io_in_0_bits_p_type),
    .io_in_0_bits_client_id(LockingRRArbiter_7_1_io_in_0_bits_client_id),
    .io_in_1_ready(LockingRRArbiter_7_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_7_1_io_in_1_valid),
    .io_in_1_bits_addr_block(LockingRRArbiter_7_1_io_in_1_bits_addr_block),
    .io_in_1_bits_p_type(LockingRRArbiter_7_1_io_in_1_bits_p_type),
    .io_in_1_bits_client_id(LockingRRArbiter_7_1_io_in_1_bits_client_id),
    .io_in_2_ready(LockingRRArbiter_7_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_7_1_io_in_2_valid),
    .io_in_2_bits_addr_block(LockingRRArbiter_7_1_io_in_2_bits_addr_block),
    .io_in_2_bits_p_type(LockingRRArbiter_7_1_io_in_2_bits_p_type),
    .io_in_2_bits_client_id(LockingRRArbiter_7_1_io_in_2_bits_client_id),
    .io_out_ready(LockingRRArbiter_7_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_7_1_io_out_valid),
    .io_out_bits_addr_block(LockingRRArbiter_7_1_io_out_bits_addr_block),
    .io_out_bits_p_type(LockingRRArbiter_7_1_io_out_bits_p_type),
    .io_out_bits_client_id(LockingRRArbiter_7_1_io_out_bits_client_id),
    .io_chosen(LockingRRArbiter_7_1_io_chosen)
  );
  LockingRRArbiter_8 LockingRRArbiter_8_1 (
    .clk(LockingRRArbiter_8_1_clk),
    .reset(LockingRRArbiter_8_1_reset),
    .io_in_0_ready(LockingRRArbiter_8_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_8_1_io_in_0_valid),
    .io_in_0_bits_addr_beat(LockingRRArbiter_8_1_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_8_1_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(LockingRRArbiter_8_1_io_in_0_bits_g_type),
    .io_in_0_bits_data(LockingRRArbiter_8_1_io_in_0_bits_data),
    .io_in_0_bits_client_id(LockingRRArbiter_8_1_io_in_0_bits_client_id),
    .io_in_1_ready(LockingRRArbiter_8_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_8_1_io_in_1_valid),
    .io_in_1_bits_addr_beat(LockingRRArbiter_8_1_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_8_1_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(LockingRRArbiter_8_1_io_in_1_bits_g_type),
    .io_in_1_bits_data(LockingRRArbiter_8_1_io_in_1_bits_data),
    .io_in_1_bits_client_id(LockingRRArbiter_8_1_io_in_1_bits_client_id),
    .io_in_2_ready(LockingRRArbiter_8_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_8_1_io_in_2_valid),
    .io_in_2_bits_addr_beat(LockingRRArbiter_8_1_io_in_2_bits_addr_beat),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_8_1_io_in_2_bits_client_xact_id),
    .io_in_2_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_g_type(LockingRRArbiter_8_1_io_in_2_bits_g_type),
    .io_in_2_bits_data(LockingRRArbiter_8_1_io_in_2_bits_data),
    .io_in_2_bits_client_id(LockingRRArbiter_8_1_io_in_2_bits_client_id),
    .io_out_ready(LockingRRArbiter_8_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_8_1_io_out_valid),
    .io_out_bits_addr_beat(LockingRRArbiter_8_1_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(LockingRRArbiter_8_1_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(LockingRRArbiter_8_1_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(LockingRRArbiter_8_1_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(LockingRRArbiter_8_1_io_out_bits_g_type),
    .io_out_bits_data(LockingRRArbiter_8_1_io_out_bits_data),
    .io_out_bits_client_id(LockingRRArbiter_8_1_io_out_bits_client_id),
    .io_chosen(LockingRRArbiter_8_1_io_chosen)
  );
  assign io_inner_acquire_ready = T_1245;
  assign io_inner_grant_valid = LockingRRArbiter_8_1_io_out_valid;
  assign io_inner_grant_bits_addr_beat = LockingRRArbiter_8_1_io_out_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = LockingRRArbiter_8_1_io_out_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = LockingRRArbiter_8_1_io_out_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = LockingRRArbiter_8_1_io_out_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = LockingRRArbiter_8_1_io_out_bits_g_type;
  assign io_inner_grant_bits_data = LockingRRArbiter_8_1_io_out_bits_data;
  assign io_inner_grant_bits_client_id = LockingRRArbiter_8_1_io_out_bits_client_id;
  assign io_inner_finish_ready = T_1324;
  assign io_inner_probe_valid = LockingRRArbiter_7_1_io_out_valid;
  assign io_inner_probe_bits_addr_block = LockingRRArbiter_7_1_io_out_bits_addr_block;
  assign io_inner_probe_bits_p_type = LockingRRArbiter_7_1_io_out_bits_p_type;
  assign io_inner_probe_bits_client_id = LockingRRArbiter_7_1_io_out_bits_client_id;
  assign io_inner_release_ready = T_1288;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_outer_acquire_bits_addr_block = outer_arb_io_out_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = outer_arb_io_out_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = outer_arb_io_out_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = outer_arb_io_out_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = outer_arb_io_out_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = outer_arb_io_out_acquire_bits_union;
  assign io_outer_acquire_bits_data = outer_arb_io_out_acquire_bits_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = outer_arb_io_out_release_valid;
  assign io_outer_release_bits_addr_beat = outer_arb_io_out_release_bits_addr_beat;
  assign io_outer_release_bits_addr_block = outer_arb_io_out_release_bits_addr_block;
  assign io_outer_release_bits_client_xact_id = outer_arb_io_out_release_bits_client_xact_id;
  assign io_outer_release_bits_voluntary = outer_arb_io_out_release_bits_voluntary;
  assign io_outer_release_bits_r_type = outer_arb_io_out_release_bits_r_type;
  assign io_outer_release_bits_data = outer_arb_io_out_release_bits_data;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = outer_arb_io_out_finish_bits_manager_xact_id;
  assign io_outer_finish_bits_manager_id = outer_arb_io_out_finish_bits_manager_id;
  assign trackerList_0_clk = clk;
  assign trackerList_0_reset = reset;
  assign trackerList_0_io_inner_acquire_valid = T_1248;
  assign trackerList_0_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign trackerList_0_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign trackerList_0_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign trackerList_0_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign trackerList_0_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign trackerList_0_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign trackerList_0_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign trackerList_0_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign trackerList_0_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_0_ready;
  assign trackerList_0_io_inner_finish_valid = T_1308;
  assign trackerList_0_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign trackerList_0_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_0_ready;
  assign trackerList_0_io_inner_release_valid = io_inner_release_valid;
  assign trackerList_0_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign trackerList_0_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign trackerList_0_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign trackerList_0_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign trackerList_0_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign trackerList_0_io_inner_release_bits_data = io_inner_release_bits_data;
  assign trackerList_0_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign trackerList_0_io_incoherent_0 = io_incoherent_0;
  assign trackerList_0_io_outer_acquire_ready = outer_arb_io_in_0_acquire_ready;
  assign trackerList_0_io_outer_probe_valid = outer_arb_io_in_0_probe_valid;
  assign trackerList_0_io_outer_probe_bits_addr_block = outer_arb_io_in_0_probe_bits_addr_block;
  assign trackerList_0_io_outer_probe_bits_p_type = outer_arb_io_in_0_probe_bits_p_type;
  assign trackerList_0_io_outer_release_ready = outer_arb_io_in_0_release_ready;
  assign trackerList_0_io_outer_grant_valid = outer_arb_io_in_0_grant_valid;
  assign trackerList_0_io_outer_grant_bits_addr_beat = outer_arb_io_in_0_grant_bits_addr_beat;
  assign trackerList_0_io_outer_grant_bits_client_xact_id = outer_arb_io_in_0_grant_bits_client_xact_id;
  assign trackerList_0_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_0_grant_bits_manager_xact_id;
  assign trackerList_0_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_0_grant_bits_is_builtin_type;
  assign trackerList_0_io_outer_grant_bits_g_type = outer_arb_io_in_0_grant_bits_g_type;
  assign trackerList_0_io_outer_grant_bits_data = outer_arb_io_in_0_grant_bits_data;
  assign trackerList_0_io_outer_grant_bits_manager_id = outer_arb_io_in_0_grant_bits_manager_id;
  assign trackerList_0_io_outer_finish_ready = outer_arb_io_in_0_finish_ready;
  assign trackerList_0_io_alloc_iacq_should = T_1251;
  assign trackerList_0_io_alloc_irel_should = T_1294;
  assign trackerList_0_io_alloc_oprb_should = GEN_0;
  assign trackerList_1_clk = clk;
  assign trackerList_1_reset = reset;
  assign trackerList_1_io_inner_acquire_valid = T_1248;
  assign trackerList_1_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign trackerList_1_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign trackerList_1_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign trackerList_1_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign trackerList_1_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign trackerList_1_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign trackerList_1_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign trackerList_1_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign trackerList_1_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_1_ready;
  assign trackerList_1_io_inner_finish_valid = T_1311;
  assign trackerList_1_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign trackerList_1_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_1_ready;
  assign trackerList_1_io_inner_release_valid = io_inner_release_valid;
  assign trackerList_1_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign trackerList_1_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign trackerList_1_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign trackerList_1_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign trackerList_1_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign trackerList_1_io_inner_release_bits_data = io_inner_release_bits_data;
  assign trackerList_1_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign trackerList_1_io_incoherent_0 = io_incoherent_0;
  assign trackerList_1_io_outer_acquire_ready = outer_arb_io_in_1_acquire_ready;
  assign trackerList_1_io_outer_probe_valid = outer_arb_io_in_1_probe_valid;
  assign trackerList_1_io_outer_probe_bits_addr_block = outer_arb_io_in_1_probe_bits_addr_block;
  assign trackerList_1_io_outer_probe_bits_p_type = outer_arb_io_in_1_probe_bits_p_type;
  assign trackerList_1_io_outer_release_ready = outer_arb_io_in_1_release_ready;
  assign trackerList_1_io_outer_grant_valid = outer_arb_io_in_1_grant_valid;
  assign trackerList_1_io_outer_grant_bits_addr_beat = outer_arb_io_in_1_grant_bits_addr_beat;
  assign trackerList_1_io_outer_grant_bits_client_xact_id = outer_arb_io_in_1_grant_bits_client_xact_id;
  assign trackerList_1_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_1_grant_bits_manager_xact_id;
  assign trackerList_1_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_1_grant_bits_is_builtin_type;
  assign trackerList_1_io_outer_grant_bits_g_type = outer_arb_io_in_1_grant_bits_g_type;
  assign trackerList_1_io_outer_grant_bits_data = outer_arb_io_in_1_grant_bits_data;
  assign trackerList_1_io_outer_grant_bits_manager_id = outer_arb_io_in_1_grant_bits_manager_id;
  assign trackerList_1_io_outer_finish_ready = outer_arb_io_in_1_finish_ready;
  assign trackerList_1_io_alloc_iacq_should = T_1256;
  assign trackerList_1_io_alloc_irel_should = T_1299;
  assign trackerList_1_io_alloc_oprb_should = GEN_1;
  assign trackerList_2_clk = clk;
  assign trackerList_2_reset = reset;
  assign trackerList_2_io_inner_acquire_valid = T_1248;
  assign trackerList_2_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign trackerList_2_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign trackerList_2_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign trackerList_2_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign trackerList_2_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign trackerList_2_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign trackerList_2_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign trackerList_2_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign trackerList_2_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_2_ready;
  assign trackerList_2_io_inner_finish_valid = T_1314;
  assign trackerList_2_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign trackerList_2_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_2_ready;
  assign trackerList_2_io_inner_release_valid = io_inner_release_valid;
  assign trackerList_2_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign trackerList_2_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign trackerList_2_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign trackerList_2_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign trackerList_2_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign trackerList_2_io_inner_release_bits_data = io_inner_release_bits_data;
  assign trackerList_2_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign trackerList_2_io_incoherent_0 = io_incoherent_0;
  assign trackerList_2_io_outer_acquire_ready = outer_arb_io_in_2_acquire_ready;
  assign trackerList_2_io_outer_probe_valid = outer_arb_io_in_2_probe_valid;
  assign trackerList_2_io_outer_probe_bits_addr_block = outer_arb_io_in_2_probe_bits_addr_block;
  assign trackerList_2_io_outer_probe_bits_p_type = outer_arb_io_in_2_probe_bits_p_type;
  assign trackerList_2_io_outer_release_ready = outer_arb_io_in_2_release_ready;
  assign trackerList_2_io_outer_grant_valid = outer_arb_io_in_2_grant_valid;
  assign trackerList_2_io_outer_grant_bits_addr_beat = outer_arb_io_in_2_grant_bits_addr_beat;
  assign trackerList_2_io_outer_grant_bits_client_xact_id = outer_arb_io_in_2_grant_bits_client_xact_id;
  assign trackerList_2_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_2_grant_bits_manager_xact_id;
  assign trackerList_2_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_2_grant_bits_is_builtin_type;
  assign trackerList_2_io_outer_grant_bits_g_type = outer_arb_io_in_2_grant_bits_g_type;
  assign trackerList_2_io_outer_grant_bits_data = outer_arb_io_in_2_grant_bits_data;
  assign trackerList_2_io_outer_grant_bits_manager_id = outer_arb_io_in_2_grant_bits_manager_id;
  assign trackerList_2_io_outer_finish_ready = outer_arb_io_in_2_finish_ready;
  assign trackerList_2_io_alloc_iacq_should = T_1261;
  assign trackerList_2_io_alloc_irel_should = T_1304;
  assign trackerList_2_io_alloc_oprb_should = GEN_2;
  assign outer_arb_clk = clk;
  assign outer_arb_reset = reset;
  assign outer_arb_io_in_0_acquire_valid = trackerList_0_io_outer_acquire_valid;
  assign outer_arb_io_in_0_acquire_bits_addr_block = trackerList_0_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_0_acquire_bits_client_xact_id = trackerList_0_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_0_acquire_bits_addr_beat = trackerList_0_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_0_acquire_bits_is_builtin_type = trackerList_0_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_0_acquire_bits_a_type = trackerList_0_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_0_acquire_bits_union = trackerList_0_io_outer_acquire_bits_union;
  assign outer_arb_io_in_0_acquire_bits_data = trackerList_0_io_outer_acquire_bits_data;
  assign outer_arb_io_in_0_probe_ready = trackerList_0_io_outer_probe_ready;
  assign outer_arb_io_in_0_release_valid = trackerList_0_io_outer_release_valid;
  assign outer_arb_io_in_0_release_bits_addr_beat = trackerList_0_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_0_release_bits_addr_block = trackerList_0_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_0_release_bits_client_xact_id = trackerList_0_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_0_release_bits_voluntary = trackerList_0_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_0_release_bits_r_type = trackerList_0_io_outer_release_bits_r_type;
  assign outer_arb_io_in_0_release_bits_data = trackerList_0_io_outer_release_bits_data;
  assign outer_arb_io_in_0_grant_ready = trackerList_0_io_outer_grant_ready;
  assign outer_arb_io_in_0_finish_valid = trackerList_0_io_outer_finish_valid;
  assign outer_arb_io_in_0_finish_bits_manager_xact_id = trackerList_0_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_0_finish_bits_manager_id = trackerList_0_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_1_acquire_valid = trackerList_1_io_outer_acquire_valid;
  assign outer_arb_io_in_1_acquire_bits_addr_block = trackerList_1_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_1_acquire_bits_client_xact_id = trackerList_1_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_1_acquire_bits_addr_beat = trackerList_1_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_1_acquire_bits_is_builtin_type = trackerList_1_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_1_acquire_bits_a_type = trackerList_1_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_1_acquire_bits_union = trackerList_1_io_outer_acquire_bits_union;
  assign outer_arb_io_in_1_acquire_bits_data = trackerList_1_io_outer_acquire_bits_data;
  assign outer_arb_io_in_1_probe_ready = trackerList_1_io_outer_probe_ready;
  assign outer_arb_io_in_1_release_valid = trackerList_1_io_outer_release_valid;
  assign outer_arb_io_in_1_release_bits_addr_beat = trackerList_1_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_1_release_bits_addr_block = trackerList_1_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_1_release_bits_client_xact_id = trackerList_1_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_1_release_bits_voluntary = trackerList_1_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_1_release_bits_r_type = trackerList_1_io_outer_release_bits_r_type;
  assign outer_arb_io_in_1_release_bits_data = trackerList_1_io_outer_release_bits_data;
  assign outer_arb_io_in_1_grant_ready = trackerList_1_io_outer_grant_ready;
  assign outer_arb_io_in_1_finish_valid = trackerList_1_io_outer_finish_valid;
  assign outer_arb_io_in_1_finish_bits_manager_xact_id = trackerList_1_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_1_finish_bits_manager_id = trackerList_1_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_2_acquire_valid = trackerList_2_io_outer_acquire_valid;
  assign outer_arb_io_in_2_acquire_bits_addr_block = trackerList_2_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_2_acquire_bits_client_xact_id = trackerList_2_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_2_acquire_bits_addr_beat = trackerList_2_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_2_acquire_bits_is_builtin_type = trackerList_2_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_2_acquire_bits_a_type = trackerList_2_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_2_acquire_bits_union = trackerList_2_io_outer_acquire_bits_union;
  assign outer_arb_io_in_2_acquire_bits_data = trackerList_2_io_outer_acquire_bits_data;
  assign outer_arb_io_in_2_probe_ready = trackerList_2_io_outer_probe_ready;
  assign outer_arb_io_in_2_release_valid = trackerList_2_io_outer_release_valid;
  assign outer_arb_io_in_2_release_bits_addr_beat = trackerList_2_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_2_release_bits_addr_block = trackerList_2_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_2_release_bits_client_xact_id = trackerList_2_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_2_release_bits_voluntary = trackerList_2_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_2_release_bits_r_type = trackerList_2_io_outer_release_bits_r_type;
  assign outer_arb_io_in_2_release_bits_data = trackerList_2_io_outer_release_bits_data;
  assign outer_arb_io_in_2_grant_ready = trackerList_2_io_outer_grant_ready;
  assign outer_arb_io_in_2_finish_valid = trackerList_2_io_outer_finish_valid;
  assign outer_arb_io_in_2_finish_bits_manager_xact_id = trackerList_2_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_2_finish_bits_manager_id = trackerList_2_io_outer_finish_bits_manager_id;
  assign outer_arb_io_out_acquire_ready = io_outer_acquire_ready;
  assign outer_arb_io_out_probe_valid = io_outer_probe_valid;
  assign outer_arb_io_out_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign outer_arb_io_out_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign outer_arb_io_out_release_ready = io_outer_release_ready;
  assign outer_arb_io_out_grant_valid = io_outer_grant_valid;
  assign outer_arb_io_out_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign outer_arb_io_out_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign outer_arb_io_out_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign outer_arb_io_out_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign outer_arb_io_out_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign outer_arb_io_out_grant_bits_data = io_outer_grant_bits_data;
  assign outer_arb_io_out_grant_bits_manager_id = io_outer_grant_bits_manager_id;
  assign outer_arb_io_out_finish_ready = io_outer_finish_ready;
  assign T_1215 = io_inner_acquire_valid & io_inner_release_valid;
  assign T_1216 = io_inner_release_bits_addr_block == io_inner_acquire_bits_addr_block;
  assign irel_vs_iacq_conflict = T_1215 & T_1216;
  assign T_1218 = irel_vs_iacq_conflict == 1'h0;
  assign T_1219 = {trackerList_2_io_inner_acquire_ready,trackerList_1_io_inner_acquire_ready};
  assign T_1220 = {T_1219,trackerList_0_io_inner_acquire_ready};
  assign T_1221 = {trackerList_2_io_alloc_iacq_can,trackerList_1_io_alloc_iacq_can};
  assign T_1222 = {T_1221,trackerList_0_io_alloc_iacq_can};
  assign T_1223 = T_1222[0];
  assign T_1224 = T_1222[1];
  assign T_1225 = T_1222[2];
  assign T_1231 = T_1225 ? 3'h4 : 3'h0;
  assign T_1232 = T_1224 ? 3'h2 : T_1231;
  assign T_1233 = T_1223 ? 3'h1 : T_1232;
  assign T_1234 = {trackerList_2_io_alloc_iacq_matches,trackerList_1_io_alloc_iacq_matches};
  assign T_1235 = {T_1234,trackerList_0_io_alloc_iacq_matches};
  assign T_1237 = T_1235 != 3'h0;
  assign T_1239 = T_1237 == 1'h0;
  assign T_1241 = T_1239 ? T_1222 : T_1235;
  assign T_1242 = T_1241 & T_1220;
  assign T_1244 = T_1242 != 3'h0;
  assign T_1245 = T_1244 & T_1218;
  assign T_1248 = io_inner_acquire_valid & T_1218;
  assign T_1249 = T_1233[0];
  assign T_1250 = T_1249 & T_1239;
  assign T_1251 = T_1250 & T_1218;
  assign T_1254 = T_1233[1];
  assign T_1255 = T_1254 & T_1239;
  assign T_1256 = T_1255 & T_1218;
  assign T_1259 = T_1233[2];
  assign T_1260 = T_1259 & T_1239;
  assign T_1261 = T_1260 & T_1218;
  assign T_1262 = {trackerList_2_io_inner_release_ready,trackerList_1_io_inner_release_ready};
  assign T_1263 = {T_1262,trackerList_0_io_inner_release_ready};
  assign T_1264 = {trackerList_2_io_alloc_irel_can,trackerList_1_io_alloc_irel_can};
  assign T_1265 = {T_1264,trackerList_0_io_alloc_irel_can};
  assign T_1266 = T_1265[0];
  assign T_1267 = T_1265[1];
  assign T_1268 = T_1265[2];
  assign T_1274 = T_1268 ? 3'h4 : 3'h0;
  assign T_1275 = T_1267 ? 3'h2 : T_1274;
  assign T_1276 = T_1266 ? 3'h1 : T_1275;
  assign T_1277 = {trackerList_2_io_alloc_irel_matches,trackerList_1_io_alloc_irel_matches};
  assign T_1278 = {T_1277,trackerList_0_io_alloc_irel_matches};
  assign T_1280 = T_1278 != 3'h0;
  assign T_1282 = T_1280 == 1'h0;
  assign T_1285 = T_1282 ? T_1265 : T_1278;
  assign T_1286 = T_1285 & T_1263;
  assign T_1288 = T_1286 != 3'h0;
  assign T_1293 = T_1276[0];
  assign T_1294 = T_1293 & T_1282;
  assign T_1298 = T_1276[1];
  assign T_1299 = T_1298 & T_1282;
  assign T_1303 = T_1276[2];
  assign T_1304 = T_1303 & T_1282;
  assign LockingRRArbiter_7_1_clk = clk;
  assign LockingRRArbiter_7_1_reset = reset;
  assign LockingRRArbiter_7_1_io_in_0_valid = trackerList_0_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_0_bits_addr_block = trackerList_0_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_0_bits_p_type = trackerList_0_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_0_bits_client_id = trackerList_0_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_1_valid = trackerList_1_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_1_bits_addr_block = trackerList_1_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_1_bits_p_type = trackerList_1_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_1_bits_client_id = trackerList_1_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_2_valid = trackerList_2_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_2_bits_addr_block = trackerList_2_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_2_bits_p_type = trackerList_2_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_2_bits_client_id = trackerList_2_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_out_ready = io_inner_probe_ready;
  assign LockingRRArbiter_8_1_clk = clk;
  assign LockingRRArbiter_8_1_reset = reset;
  assign LockingRRArbiter_8_1_io_in_0_valid = trackerList_0_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_0_bits_addr_beat = trackerList_0_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_0_bits_client_xact_id = trackerList_0_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_0_bits_manager_xact_id = trackerList_0_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_0_bits_is_builtin_type = trackerList_0_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_0_bits_g_type = trackerList_0_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_0_bits_data = trackerList_0_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_0_bits_client_id = trackerList_0_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_1_valid = trackerList_1_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_1_bits_addr_beat = trackerList_1_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_1_bits_client_xact_id = trackerList_1_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_1_bits_manager_xact_id = trackerList_1_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_1_bits_is_builtin_type = trackerList_1_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_1_bits_g_type = trackerList_1_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_1_bits_data = trackerList_1_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_1_bits_client_id = trackerList_1_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_2_valid = trackerList_2_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_2_bits_addr_beat = trackerList_2_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_2_bits_client_xact_id = trackerList_2_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_2_bits_manager_xact_id = trackerList_2_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_2_bits_is_builtin_type = trackerList_2_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_2_bits_g_type = trackerList_2_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_2_bits_data = trackerList_2_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_2_bits_client_id = trackerList_2_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_out_ready = io_inner_grant_ready;
  assign T_1307 = io_inner_finish_bits_manager_xact_id == 2'h0;
  assign T_1308 = io_inner_finish_valid & T_1307;
  assign T_1310 = io_inner_finish_bits_manager_xact_id == 2'h1;
  assign T_1311 = io_inner_finish_valid & T_1310;
  assign T_1313 = io_inner_finish_bits_manager_xact_id == 2'h2;
  assign T_1314 = io_inner_finish_valid & T_1313;
  assign T_1316 = io_inner_finish_bits_manager_xact_id & 2'h1;
  assign T_1318 = io_inner_finish_bits_manager_xact_id >= 2'h2;
  assign T_1322 = T_1316 >= 2'h1;
  assign T_1323 = T_1322 ? trackerList_1_io_inner_finish_ready : trackerList_0_io_inner_finish_ready;
  assign T_1324 = T_1318 ? trackerList_2_io_inner_finish_ready : T_1323;
  assign T_1328 = io_outer_probe_valid == 1'h0;
  assign T_1329 = T_1328 | reset;
  assign T_1331 = T_1329 == 1'h0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_0 = GEN_3[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_4[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_5[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_3 = {1{$random}};
  GEN_4 = {1{$random}};
  GEN_5 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1331) begin
          $fwrite(32'h80000002,"Assertion failed: L2 agent got illegal probe\n    at Agents.scala:160 assert(!io.outer.probe.valid, \"L2 agent got illegal probe\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1331) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module MMIOTileLinkManager(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input   io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output  io_inner_grant_bits_client_xact_id,
  output [1:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [1:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input   io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data
);
  wire  T_880;
  wire [2:0] T_889_0;
  wire  T_891;
  wire  T_892;
  wire  multibeat_fire;
  wire  T_894;
  wire  multibeat_start;
  wire  T_896;
  wire  multibeat_end;
  reg [3:0] xact_pending;
  reg [31:0] GEN_31;
  wire [3:0] T_898;
  wire  T_899;
  wire  T_900;
  wire  T_901;
  wire [1:0] T_907;
  wire [1:0] T_908;
  wire [1:0] xact_id_sel;
  reg [1:0] xact_id_reg;
  reg [31:0] GEN_32;
  wire [1:0] GEN_4;
  reg  xact_multibeat;
  reg [31:0] GEN_33;
  wire [1:0] outer_xact_id;
  wire  T_912;
  wire  xact_free;
  reg  xact_buffer_0_client_id;
  reg [31:0] GEN_34;
  reg  xact_buffer_0_client_xact_id;
  reg [31:0] GEN_35;
  reg  xact_buffer_1_client_id;
  reg [31:0] GEN_36;
  reg  xact_buffer_1_client_xact_id;
  reg [31:0] GEN_37;
  reg  xact_buffer_2_client_id;
  reg [31:0] GEN_38;
  reg  xact_buffer_2_client_xact_id;
  reg [31:0] GEN_39;
  reg  xact_buffer_3_client_id;
  reg [31:0] GEN_40;
  reg  xact_buffer_3_client_xact_id;
  reg [31:0] GEN_41;
  wire  T_1229;
  wire  T_1230;
  wire [2:0] T_1240_0;
  wire  T_1242;
  wire  T_1243;
  wire  T_1245;
  wire  T_1248;
  wire  T_1249;
  wire [3:0] T_1251;
  wire [3:0] T_1253;
  wire [3:0] T_1254;
  wire  T_1255;
  wire [3:0] T_1257;
  wire [3:0] T_1259;
  wire [3:0] T_1260;
  wire [3:0] T_1261;
  wire  T_1262;
  wire [2:0] T_1270_0;
  wire [3:0] GEN_2;
  wire  T_1272;
  wire  T_1273;
  wire  T_1274;
  wire  T_1277;
  wire  T_1279;
  wire  T_1280;
  wire  T_1281;
  wire  T_1287;
  wire  T_1289;
  wire  T_1292;
  wire  T_1293;
  wire [3:0] T_1295;
  wire [3:0] T_1297;
  wire [3:0] T_1298;
  wire [3:0] T_1299;
  wire [2:0] T_1309_0;
  wire  T_1311;
  wire  T_1312;
  wire  T_1314;
  wire  T_1317;
  wire  T_1318;
  wire  GEN_0;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_1;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_2_client_id;
  wire  GEN_2_client_xact_id;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_3_client_id;
  wire  GEN_3_client_xact_id;
  wire [25:0] GEN_3;
  reg [31:0] GEN_42;
  wire [1:0] GEN_13;
  reg [31:0] GEN_43;
  wire  GEN_18;
  reg [31:0] GEN_44;
  assign io_inner_acquire_ready = T_1229;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = GEN_3_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_client_id = GEN_2_client_id;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_3;
  assign io_inner_probe_bits_p_type = GEN_13;
  assign io_inner_probe_bits_client_id = GEN_18;
  assign io_inner_release_ready = 1'h0;
  assign io_outer_acquire_valid = T_1230;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = outer_xact_id;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign T_880 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_889_0 = 3'h3;
  assign T_891 = io_outer_acquire_bits_a_type == T_889_0;
  assign T_892 = io_outer_acquire_bits_is_builtin_type & T_891;
  assign multibeat_fire = T_880 & T_892;
  assign T_894 = io_outer_acquire_bits_addr_beat == 3'h0;
  assign multibeat_start = multibeat_fire & T_894;
  assign T_896 = io_outer_acquire_bits_addr_beat == 3'h7;
  assign multibeat_end = multibeat_fire & T_896;
  assign T_898 = ~ xact_pending;
  assign T_899 = T_898[0];
  assign T_900 = T_898[1];
  assign T_901 = T_898[2];
  assign T_907 = T_901 ? 2'h2 : 2'h3;
  assign T_908 = T_900 ? 2'h1 : T_907;
  assign xact_id_sel = T_899 ? 2'h0 : T_908;
  assign GEN_4 = multibeat_start ? xact_id_sel : xact_id_reg;
  assign outer_xact_id = xact_multibeat ? xact_id_reg : xact_id_sel;
  assign T_912 = T_898 == 4'h0;
  assign xact_free = T_912 == 1'h0;
  assign T_1229 = io_outer_acquire_ready & xact_free;
  assign T_1230 = io_inner_acquire_valid & xact_free;
  assign T_1240_0 = 3'h3;
  assign T_1242 = io_outer_acquire_bits_a_type == T_1240_0;
  assign T_1243 = io_outer_acquire_bits_is_builtin_type & T_1242;
  assign T_1245 = T_1243 == 1'h0;
  assign T_1248 = T_1245 | T_896;
  assign T_1249 = T_880 & T_1248;
  assign T_1251 = 4'h1 << io_outer_acquire_bits_client_xact_id;
  assign T_1253 = T_1249 ? T_1251 : 4'h0;
  assign T_1254 = xact_pending | T_1253;
  assign T_1255 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_1257 = 4'h1 << io_inner_finish_bits_manager_xact_id;
  assign T_1259 = T_1255 ? T_1257 : 4'h0;
  assign T_1260 = ~ T_1259;
  assign T_1261 = T_1254 & T_1260;
  assign T_1262 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_1270_0 = 3'h5;
  assign GEN_2 = {{1'd0}, T_1270_0};
  assign T_1272 = io_inner_grant_bits_g_type == GEN_2;
  assign T_1273 = io_inner_grant_bits_g_type == 4'h0;
  assign T_1274 = io_inner_grant_bits_is_builtin_type ? T_1272 : T_1273;
  assign T_1277 = T_1274 == 1'h0;
  assign T_1279 = io_inner_grant_bits_addr_beat == 3'h7;
  assign T_1280 = T_1277 | T_1279;
  assign T_1281 = T_1262 & T_1280;
  assign T_1287 = io_inner_grant_bits_is_builtin_type & T_1273;
  assign T_1289 = T_1287 == 1'h0;
  assign T_1292 = T_1289 == 1'h0;
  assign T_1293 = T_1281 & T_1292;
  assign T_1295 = 4'h1 << io_inner_grant_bits_manager_xact_id;
  assign T_1297 = T_1293 ? T_1295 : 4'h0;
  assign T_1298 = ~ T_1297;
  assign T_1299 = T_1261 & T_1298;
  assign T_1309_0 = 3'h3;
  assign T_1311 = io_outer_acquire_bits_a_type == T_1309_0;
  assign T_1312 = io_outer_acquire_bits_is_builtin_type & T_1311;
  assign T_1314 = T_1312 == 1'h0;
  assign T_1317 = T_1314 | T_896;
  assign T_1318 = T_880 & T_1317;
  assign GEN_0 = io_inner_acquire_bits_client_id;
  assign GEN_5 = 2'h0 == outer_xact_id ? GEN_0 : xact_buffer_0_client_id;
  assign GEN_6 = 2'h1 == outer_xact_id ? GEN_0 : xact_buffer_1_client_id;
  assign GEN_7 = 2'h2 == outer_xact_id ? GEN_0 : xact_buffer_2_client_id;
  assign GEN_8 = 2'h3 == outer_xact_id ? GEN_0 : xact_buffer_3_client_id;
  assign GEN_1 = io_inner_acquire_bits_client_xact_id;
  assign GEN_9 = 2'h0 == outer_xact_id ? GEN_1 : xact_buffer_0_client_xact_id;
  assign GEN_10 = 2'h1 == outer_xact_id ? GEN_1 : xact_buffer_1_client_xact_id;
  assign GEN_11 = 2'h2 == outer_xact_id ? GEN_1 : xact_buffer_2_client_xact_id;
  assign GEN_12 = 2'h3 == outer_xact_id ? GEN_1 : xact_buffer_3_client_xact_id;
  assign GEN_14 = T_1318 ? GEN_5 : xact_buffer_0_client_id;
  assign GEN_15 = T_1318 ? GEN_6 : xact_buffer_1_client_id;
  assign GEN_16 = T_1318 ? GEN_7 : xact_buffer_2_client_id;
  assign GEN_17 = T_1318 ? GEN_8 : xact_buffer_3_client_id;
  assign GEN_19 = T_1318 ? GEN_9 : xact_buffer_0_client_xact_id;
  assign GEN_20 = T_1318 ? GEN_10 : xact_buffer_1_client_xact_id;
  assign GEN_21 = T_1318 ? GEN_11 : xact_buffer_2_client_xact_id;
  assign GEN_22 = T_1318 ? GEN_12 : xact_buffer_3_client_xact_id;
  assign GEN_23 = multibeat_start ? 1'h1 : xact_multibeat;
  assign GEN_24 = multibeat_end ? 1'h0 : GEN_23;
  assign GEN_2_client_id = GEN_29;
  assign GEN_2_client_xact_id = GEN_30;
  assign GEN_25 = 2'h1 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_id : xact_buffer_0_client_id;
  assign GEN_26 = 2'h1 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_xact_id : xact_buffer_0_client_xact_id;
  assign GEN_27 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_id : GEN_25;
  assign GEN_28 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_xact_id : GEN_26;
  assign GEN_29 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_id : GEN_27;
  assign GEN_30 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_xact_id : GEN_28;
  assign GEN_3_client_id = GEN_29;
  assign GEN_3_client_xact_id = GEN_30;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_42[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_13 = GEN_43[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_18 = GEN_44[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  xact_pending = GEN_31[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  xact_id_reg = GEN_32[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  xact_multibeat = GEN_33[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  xact_buffer_0_client_id = GEN_34[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {1{$random}};
  xact_buffer_0_client_xact_id = GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  xact_buffer_1_client_id = GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  xact_buffer_1_client_xact_id = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {1{$random}};
  xact_buffer_2_client_id = GEN_38[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  xact_buffer_2_client_xact_id = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  xact_buffer_3_client_id = GEN_40[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  xact_buffer_3_client_xact_id = GEN_41[0:0];
  `endif
  GEN_42 = {1{$random}};
  GEN_43 = {1{$random}};
  GEN_44 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      xact_pending <= 4'h0;
    end else begin
      xact_pending <= T_1299;
    end
    if(1'h0) begin
    end else begin
      if(multibeat_start) begin
        if(T_899) begin
          xact_id_reg <= 2'h0;
        end else begin
          if(T_900) begin
            xact_id_reg <= 2'h1;
          end else begin
            if(T_901) begin
              xact_id_reg <= 2'h2;
            end else begin
              xact_id_reg <= 2'h3;
            end
          end
        end
      end
    end
    if(reset) begin
      xact_multibeat <= 1'h0;
    end else begin
      if(multibeat_end) begin
        xact_multibeat <= 1'h0;
      end else begin
        if(multibeat_start) begin
          xact_multibeat <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h0 == outer_xact_id) begin
          xact_buffer_0_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h0 == outer_xact_id) begin
          xact_buffer_0_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h1 == outer_xact_id) begin
          xact_buffer_1_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h1 == outer_xact_id) begin
          xact_buffer_1_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h2 == outer_xact_id) begin
          xact_buffer_2_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h2 == outer_xact_id) begin
          xact_buffer_2_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h3 == outer_xact_id) begin
          xact_buffer_3_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h3 == outer_xact_id) begin
          xact_buffer_3_client_xact_id <= GEN_1;
        end
      end
    end
  end
endmodule
module ClientUncachedTileLinkIOArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [1:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [10:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [1:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module TileLinkMemoryInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data
);
  wire  ClientUncachedTileLinkIOArbiter_1_1_clk;
  wire  ClientUncachedTileLinkIOArbiter_1_1_reset;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data;
  wire [25:0] T_3009;
  ClientUncachedTileLinkIOArbiter_1 ClientUncachedTileLinkIOArbiter_1_1 (
    .clk(ClientUncachedTileLinkIOArbiter_1_1_clk),
    .reset(ClientUncachedTileLinkIOArbiter_1_1_reset),
    .io_in_0_acquire_ready(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data),
    .io_out_acquire_ready(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready),
    .io_out_acquire_valid(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready),
    .io_out_grant_valid(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = T_3009;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_clk = clk;
  assign ClientUncachedTileLinkIOArbiter_1_1_reset = reset;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data = io_out_0_grant_bits_data;
  assign T_3009 = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block >> 1'h0;
endmodule
module LockingRRArbiter_9(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [10:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [10:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [10:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [25:0] GEN_0_bits_addr_block;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire [2:0] GEN_0_bits_addr_beat;
  wire  GEN_0_bits_is_builtin_type;
  wire [2:0] GEN_0_bits_a_type;
  wire [10:0] GEN_0_bits_union;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_8;
  wire  GEN_9;
  wire [25:0] GEN_10;
  wire [1:0] GEN_11;
  wire [2:0] GEN_12;
  wire  GEN_13;
  wire [2:0] GEN_14;
  wire [10:0] GEN_15;
  wire [63:0] GEN_16;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [25:0] GEN_1_bits_addr_block;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire [2:0] GEN_1_bits_addr_beat;
  wire  GEN_1_bits_is_builtin_type;
  wire [2:0] GEN_1_bits_a_type;
  wire [10:0] GEN_1_bits_union;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [25:0] GEN_2_bits_addr_block;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire [2:0] GEN_2_bits_addr_beat;
  wire  GEN_2_bits_is_builtin_type;
  wire [2:0] GEN_2_bits_a_type;
  wire [10:0] GEN_2_bits_union;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [25:0] GEN_3_bits_addr_block;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire [2:0] GEN_3_bits_addr_beat;
  wire  GEN_3_bits_is_builtin_type;
  wire [2:0] GEN_3_bits_a_type;
  wire [10:0] GEN_3_bits_union;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [25:0] GEN_4_bits_addr_block;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire [2:0] GEN_4_bits_addr_beat;
  wire  GEN_4_bits_is_builtin_type;
  wire [2:0] GEN_4_bits_a_type;
  wire [10:0] GEN_4_bits_union;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [25:0] GEN_5_bits_addr_block;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire [2:0] GEN_5_bits_addr_beat;
  wire  GEN_5_bits_is_builtin_type;
  wire [2:0] GEN_5_bits_a_type;
  wire [10:0] GEN_5_bits_union;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [25:0] GEN_6_bits_addr_block;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire [2:0] GEN_6_bits_addr_beat;
  wire  GEN_6_bits_is_builtin_type;
  wire [2:0] GEN_6_bits_a_type;
  wire [10:0] GEN_6_bits_union;
  wire [63:0] GEN_6_bits_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [25:0] GEN_7_bits_addr_block;
  wire [1:0] GEN_7_bits_client_xact_id;
  wire [2:0] GEN_7_bits_addr_beat;
  wire  GEN_7_bits_is_builtin_type;
  wire [2:0] GEN_7_bits_a_type;
  wire [10:0] GEN_7_bits_union;
  wire [63:0] GEN_7_bits_data;
  reg [2:0] T_766;
  reg [31:0] GEN_0;
  reg  T_768;
  reg [31:0] GEN_1;
  wire  T_770;
  wire [2:0] T_779_0;
  wire  T_781;
  wire  T_782;
  wire  T_783;
  wire  T_784;
  wire [3:0] T_788;
  wire [2:0] T_789;
  wire  GEN_80;
  wire [2:0] GEN_81;
  wire  GEN_82;
  reg  lastGrant;
  reg [31:0] GEN_2;
  wire  GEN_83;
  wire  grantMask_1;
  wire  validMask_1;
  wire  T_795;
  wire  T_799;
  wire  T_801;
  wire  T_805;
  wire  T_807;
  wire  T_808;
  wire  T_809;
  wire  T_812;
  wire  T_813;
  wire  GEN_84;
  wire  GEN_85;
  assign io_in_0_ready = T_809;
  assign io_in_1_ready = T_813;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_block = GEN_1_bits_addr_block;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_addr_beat = GEN_3_bits_addr_beat;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_a_type = GEN_5_bits_a_type;
  assign io_out_bits_union = GEN_6_bits_union;
  assign io_out_bits_data = GEN_7_bits_data;
  assign io_chosen = GEN_82;
  assign choice = GEN_85;
  assign GEN_0_ready = GEN_8;
  assign GEN_0_valid = GEN_9;
  assign GEN_0_bits_addr_block = GEN_10;
  assign GEN_0_bits_client_xact_id = GEN_11;
  assign GEN_0_bits_addr_beat = GEN_12;
  assign GEN_0_bits_is_builtin_type = GEN_13;
  assign GEN_0_bits_a_type = GEN_14;
  assign GEN_0_bits_union = GEN_15;
  assign GEN_0_bits_data = GEN_16;
  assign GEN_8 = io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_9 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_13 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_14 = io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_15 = io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_16 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_1_ready = GEN_8;
  assign GEN_1_valid = GEN_9;
  assign GEN_1_bits_addr_block = GEN_10;
  assign GEN_1_bits_client_xact_id = GEN_11;
  assign GEN_1_bits_addr_beat = GEN_12;
  assign GEN_1_bits_is_builtin_type = GEN_13;
  assign GEN_1_bits_a_type = GEN_14;
  assign GEN_1_bits_union = GEN_15;
  assign GEN_1_bits_data = GEN_16;
  assign GEN_2_ready = GEN_8;
  assign GEN_2_valid = GEN_9;
  assign GEN_2_bits_addr_block = GEN_10;
  assign GEN_2_bits_client_xact_id = GEN_11;
  assign GEN_2_bits_addr_beat = GEN_12;
  assign GEN_2_bits_is_builtin_type = GEN_13;
  assign GEN_2_bits_a_type = GEN_14;
  assign GEN_2_bits_union = GEN_15;
  assign GEN_2_bits_data = GEN_16;
  assign GEN_3_ready = GEN_8;
  assign GEN_3_valid = GEN_9;
  assign GEN_3_bits_addr_block = GEN_10;
  assign GEN_3_bits_client_xact_id = GEN_11;
  assign GEN_3_bits_addr_beat = GEN_12;
  assign GEN_3_bits_is_builtin_type = GEN_13;
  assign GEN_3_bits_a_type = GEN_14;
  assign GEN_3_bits_union = GEN_15;
  assign GEN_3_bits_data = GEN_16;
  assign GEN_4_ready = GEN_8;
  assign GEN_4_valid = GEN_9;
  assign GEN_4_bits_addr_block = GEN_10;
  assign GEN_4_bits_client_xact_id = GEN_11;
  assign GEN_4_bits_addr_beat = GEN_12;
  assign GEN_4_bits_is_builtin_type = GEN_13;
  assign GEN_4_bits_a_type = GEN_14;
  assign GEN_4_bits_union = GEN_15;
  assign GEN_4_bits_data = GEN_16;
  assign GEN_5_ready = GEN_8;
  assign GEN_5_valid = GEN_9;
  assign GEN_5_bits_addr_block = GEN_10;
  assign GEN_5_bits_client_xact_id = GEN_11;
  assign GEN_5_bits_addr_beat = GEN_12;
  assign GEN_5_bits_is_builtin_type = GEN_13;
  assign GEN_5_bits_a_type = GEN_14;
  assign GEN_5_bits_union = GEN_15;
  assign GEN_5_bits_data = GEN_16;
  assign GEN_6_ready = GEN_8;
  assign GEN_6_valid = GEN_9;
  assign GEN_6_bits_addr_block = GEN_10;
  assign GEN_6_bits_client_xact_id = GEN_11;
  assign GEN_6_bits_addr_beat = GEN_12;
  assign GEN_6_bits_is_builtin_type = GEN_13;
  assign GEN_6_bits_a_type = GEN_14;
  assign GEN_6_bits_union = GEN_15;
  assign GEN_6_bits_data = GEN_16;
  assign GEN_7_ready = GEN_8;
  assign GEN_7_valid = GEN_9;
  assign GEN_7_bits_addr_block = GEN_10;
  assign GEN_7_bits_client_xact_id = GEN_11;
  assign GEN_7_bits_addr_beat = GEN_12;
  assign GEN_7_bits_is_builtin_type = GEN_13;
  assign GEN_7_bits_a_type = GEN_14;
  assign GEN_7_bits_union = GEN_15;
  assign GEN_7_bits_data = GEN_16;
  assign T_770 = T_766 != 3'h0;
  assign T_779_0 = 3'h3;
  assign T_781 = io_out_bits_a_type == T_779_0;
  assign T_782 = io_out_bits_is_builtin_type & T_781;
  assign T_783 = io_out_ready & io_out_valid;
  assign T_784 = T_783 & T_782;
  assign T_788 = T_766 + 3'h1;
  assign T_789 = T_788[2:0];
  assign GEN_80 = T_784 ? io_chosen : T_768;
  assign GEN_81 = T_784 ? T_789 : T_766;
  assign GEN_82 = T_770 ? T_768 : choice;
  assign GEN_83 = T_783 ? io_chosen : lastGrant;
  assign grantMask_1 = 1'h1 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign T_795 = validMask_1 | io_in_0_valid;
  assign T_799 = validMask_1 == 1'h0;
  assign T_801 = T_795 == 1'h0;
  assign T_805 = grantMask_1 | T_801;
  assign T_807 = T_768 == 1'h0;
  assign T_808 = T_770 ? T_807 : T_799;
  assign T_809 = T_808 & io_out_ready;
  assign T_812 = T_770 ? T_768 : T_805;
  assign T_813 = T_812 & io_out_ready;
  assign GEN_84 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_85 = validMask_1 ? 1'h1 : GEN_84;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_766 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_768 = GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_766 <= 3'h0;
    end else begin
      if(T_784) begin
        T_766 <= T_789;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_784) begin
        T_768 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_783) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ReorderQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_data,
  input  [1:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [1:0] io_deq_tag,
  output  io_deq_data,
  output  io_deq_matches
);
  reg  T_31 [0:3];
  reg [31:0] GEN_14;
  wire  T_31_T_47_data;
  wire [1:0] T_31_T_47_addr;
  wire  T_31_T_47_en;
  wire  T_31_T_51_data;
  wire [1:0] T_31_T_51_addr;
  wire  T_31_T_51_mask;
  wire  T_31_T_51_en;
  wire  T_41_0;
  wire  T_41_1;
  wire  T_41_2;
  wire  T_41_3;
  reg  T_45_0;
  reg [31:0] GEN_15;
  reg  T_45_1;
  reg [31:0] GEN_16;
  reg  T_45_2;
  reg [31:0] GEN_17;
  reg  T_45_3;
  reg [31:0] GEN_18;
  wire  GEN_0;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_1;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  T_49;
  wire  T_50;
  wire  GEN_2;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_3;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  assign io_enq_ready = GEN_0;
  assign io_deq_data = T_31_T_47_data;
  assign io_deq_matches = T_49;
  assign T_31_T_47_addr = io_deq_tag;
  assign T_31_T_47_en = 1'h1;
  assign T_31_T_47_data = T_31[T_31_T_47_addr];
  assign T_31_T_51_data = io_enq_bits_data;
  assign T_31_T_51_addr = io_enq_bits_tag;
  assign T_31_T_51_mask = T_50;
  assign T_31_T_51_en = T_50;
  assign T_41_0 = 1'h1;
  assign T_41_1 = 1'h1;
  assign T_41_2 = 1'h1;
  assign T_41_3 = 1'h1;
  assign GEN_0 = GEN_6;
  assign GEN_4 = 2'h1 == io_enq_bits_tag ? T_45_1 : T_45_0;
  assign GEN_5 = 2'h2 == io_enq_bits_tag ? T_45_2 : GEN_4;
  assign GEN_6 = 2'h3 == io_enq_bits_tag ? T_45_3 : GEN_5;
  assign GEN_1 = GEN_9;
  assign GEN_7 = 2'h1 == io_deq_tag ? T_45_1 : T_45_0;
  assign GEN_8 = 2'h2 == io_deq_tag ? T_45_2 : GEN_7;
  assign GEN_9 = 2'h3 == io_deq_tag ? T_45_3 : GEN_8;
  assign T_49 = GEN_1 == 1'h0;
  assign T_50 = io_enq_valid & io_enq_ready;
  assign GEN_2 = 1'h0;
  assign GEN_10 = 2'h0 == io_enq_bits_tag ? GEN_2 : T_45_0;
  assign GEN_11 = 2'h1 == io_enq_bits_tag ? GEN_2 : T_45_1;
  assign GEN_12 = 2'h2 == io_enq_bits_tag ? GEN_2 : T_45_2;
  assign GEN_13 = 2'h3 == io_enq_bits_tag ? GEN_2 : T_45_3;
  assign GEN_20 = T_50 ? GEN_10 : T_45_0;
  assign GEN_21 = T_50 ? GEN_11 : T_45_1;
  assign GEN_22 = T_50 ? GEN_12 : T_45_2;
  assign GEN_23 = T_50 ? GEN_13 : T_45_3;
  assign GEN_3 = 1'h1;
  assign GEN_24 = 2'h0 == io_deq_tag ? GEN_3 : GEN_20;
  assign GEN_25 = 2'h1 == io_deq_tag ? GEN_3 : GEN_21;
  assign GEN_26 = 2'h2 == io_deq_tag ? GEN_3 : GEN_22;
  assign GEN_27 = 2'h3 == io_deq_tag ? GEN_3 : GEN_23;
  assign GEN_29 = io_deq_valid ? GEN_24 : GEN_20;
  assign GEN_30 = io_deq_valid ? GEN_25 : GEN_21;
  assign GEN_31 = io_deq_valid ? GEN_26 : GEN_22;
  assign GEN_32 = io_deq_valid ? GEN_27 : GEN_23;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_14 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    T_31[initvar] = GEN_14[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_15 = {1{$random}};
  T_45_0 = GEN_15[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_16 = {1{$random}};
  T_45_1 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {1{$random}};
  T_45_2 = GEN_17[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {1{$random}};
  T_45_3 = GEN_18[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(T_31_T_51_en & T_31_T_51_mask) begin
      T_31[T_31_T_51_addr] <= T_31_T_51_data;
    end
    if(reset) begin
      T_45_0 <= T_41_0;
    end else begin
      if(io_deq_valid) begin
        if(2'h0 == io_deq_tag) begin
          T_45_0 <= GEN_3;
        end else begin
          if(T_50) begin
            if(2'h0 == io_enq_bits_tag) begin
              T_45_0 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_50) begin
          if(2'h0 == io_enq_bits_tag) begin
            T_45_0 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_45_1 <= T_41_1;
    end else begin
      if(io_deq_valid) begin
        if(2'h1 == io_deq_tag) begin
          T_45_1 <= GEN_3;
        end else begin
          if(T_50) begin
            if(2'h1 == io_enq_bits_tag) begin
              T_45_1 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_50) begin
          if(2'h1 == io_enq_bits_tag) begin
            T_45_1 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_45_2 <= T_41_2;
    end else begin
      if(io_deq_valid) begin
        if(2'h2 == io_deq_tag) begin
          T_45_2 <= GEN_3;
        end else begin
          if(T_50) begin
            if(2'h2 == io_enq_bits_tag) begin
              T_45_2 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_50) begin
          if(2'h2 == io_enq_bits_tag) begin
            T_45_2 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_45_3 <= T_41_3;
    end else begin
      if(io_deq_valid) begin
        if(2'h3 == io_deq_tag) begin
          T_45_3 <= GEN_3;
        end else begin
          if(T_50) begin
            if(2'h3 == io_enq_bits_tag) begin
              T_45_3 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_50) begin
          if(2'h3 == io_enq_bits_tag) begin
            T_45_3 <= GEN_2;
          end
        end
      end
    end
  end
endmodule
module ClientTileLinkIOUnwrapper(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [10:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_probe_ready,
  output  io_in_probe_valid,
  output [25:0] io_in_probe_bits_addr_block,
  output [1:0] io_in_probe_bits_p_type,
  output  io_in_release_ready,
  input   io_in_release_valid,
  input  [2:0] io_in_release_bits_addr_beat,
  input  [25:0] io_in_release_bits_addr_block,
  input  [1:0] io_in_release_bits_client_xact_id,
  input   io_in_release_bits_voluntary,
  input  [2:0] io_in_release_bits_r_type,
  input  [63:0] io_in_release_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  output  io_in_grant_bits_manager_id,
  output  io_in_finish_ready,
  input   io_in_finish_valid,
  input   io_in_finish_bits_manager_xact_id,
  input   io_in_finish_bits_manager_id,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [1:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [10:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [1:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  wire  acqArb_clk;
  wire  acqArb_reset;
  wire  acqArb_io_in_0_ready;
  wire  acqArb_io_in_0_valid;
  wire [25:0] acqArb_io_in_0_bits_addr_block;
  wire [1:0] acqArb_io_in_0_bits_client_xact_id;
  wire [2:0] acqArb_io_in_0_bits_addr_beat;
  wire  acqArb_io_in_0_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_0_bits_a_type;
  wire [10:0] acqArb_io_in_0_bits_union;
  wire [63:0] acqArb_io_in_0_bits_data;
  wire  acqArb_io_in_1_ready;
  wire  acqArb_io_in_1_valid;
  wire [25:0] acqArb_io_in_1_bits_addr_block;
  wire [1:0] acqArb_io_in_1_bits_client_xact_id;
  wire [2:0] acqArb_io_in_1_bits_addr_beat;
  wire  acqArb_io_in_1_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_1_bits_a_type;
  wire [10:0] acqArb_io_in_1_bits_union;
  wire [63:0] acqArb_io_in_1_bits_data;
  wire  acqArb_io_out_ready;
  wire  acqArb_io_out_valid;
  wire [25:0] acqArb_io_out_bits_addr_block;
  wire [1:0] acqArb_io_out_bits_client_xact_id;
  wire [2:0] acqArb_io_out_bits_addr_beat;
  wire  acqArb_io_out_bits_is_builtin_type;
  wire [2:0] acqArb_io_out_bits_a_type;
  wire [10:0] acqArb_io_out_bits_union;
  wire [63:0] acqArb_io_out_bits_data;
  wire  acqArb_io_chosen;
  wire  acqRoq_clk;
  wire  acqRoq_reset;
  wire  acqRoq_io_enq_ready;
  wire  acqRoq_io_enq_valid;
  wire  acqRoq_io_enq_bits_data;
  wire [1:0] acqRoq_io_enq_bits_tag;
  wire  acqRoq_io_deq_valid;
  wire [1:0] acqRoq_io_deq_tag;
  wire  acqRoq_io_deq_data;
  wire  acqRoq_io_deq_matches;
  wire  relRoq_clk;
  wire  relRoq_reset;
  wire  relRoq_io_enq_ready;
  wire  relRoq_io_enq_valid;
  wire  relRoq_io_enq_bits_data;
  wire [1:0] relRoq_io_enq_bits_tag;
  wire  relRoq_io_deq_valid;
  wire [1:0] relRoq_io_deq_tag;
  wire  relRoq_io_deq_data;
  wire  relRoq_io_deq_matches;
  wire [2:0] T_1366_0;
  wire  T_1368;
  wire  T_1369;
  wire  T_1371;
  wire  T_1373;
  wire  acq_roq_enq;
  wire  T_1375;
  wire  T_1376;
  wire  T_1377;
  wire  T_1378;
  wire  T_1379;
  wire  T_1382;
  wire  T_1384;
  wire  rel_roq_enq;
  wire  T_1386;
  wire  acq_roq_ready;
  wire  T_1388;
  wire  rel_roq_ready;
  wire  T_1389;
  wire  T_1390;
  wire  T_1391;
  wire [2:0] T_1394;
  wire [25:0] T_1423_addr_block;
  wire [1:0] T_1423_client_xact_id;
  wire [2:0] T_1423_addr_beat;
  wire  T_1423_is_builtin_type;
  wire [2:0] T_1423_a_type;
  wire [10:0] T_1423_union;
  wire [63:0] T_1423_data;
  wire  T_1451;
  wire  T_1452;
  wire  T_1453;
  wire  T_1454;
  wire [25:0] T_1577_addr_block;
  wire [1:0] T_1577_client_xact_id;
  wire [2:0] T_1577_addr_beat;
  wire  T_1577_is_builtin_type;
  wire [2:0] T_1577_a_type;
  wire [10:0] T_1577_union;
  wire [63:0] T_1577_data;
  wire  T_1605;
  wire  T_1606;
  wire [2:0] T_1614_0;
  wire [3:0] GEN_0;
  wire  T_1616;
  wire  T_1617;
  wire  T_1618;
  wire  T_1621;
  wire  T_1623;
  wire  T_1624;
  wire  grant_deq_roq;
  wire  T_1625;
  wire  T_1627;
  wire  T_1628;
  wire  T_1630;
  wire  T_1631;
  wire  T_1632;
  wire  T_1633;
  wire  T_1635;
  wire [3:0] T_1636;
  wire [2:0] acq_grant_addr_beat;
  wire [1:0] acq_grant_client_xact_id;
  wire  acq_grant_manager_xact_id;
  wire  acq_grant_is_builtin_type;
  wire [3:0] acq_grant_g_type;
  wire [63:0] acq_grant_data;
  wire  T_1691;
  wire  T_1692;
  wire  T_1693;
  wire  T_1695;
  wire [2:0] rel_grant_addr_beat;
  wire [1:0] rel_grant_client_xact_id;
  wire  rel_grant_manager_xact_id;
  wire  rel_grant_is_builtin_type;
  wire [3:0] rel_grant_g_type;
  wire [63:0] rel_grant_data;
  wire [2:0] T_1751_addr_beat;
  wire [1:0] T_1751_client_xact_id;
  wire  T_1751_manager_xact_id;
  wire  T_1751_is_builtin_type;
  wire [3:0] T_1751_g_type;
  wire [63:0] T_1751_data;
  wire [25:0] GEN_1;
  reg [31:0] GEN_4;
  wire [1:0] GEN_2;
  reg [31:0] GEN_5;
  wire  GEN_3;
  reg [31:0] GEN_6;
  LockingRRArbiter_9 acqArb (
    .clk(acqArb_clk),
    .reset(acqArb_reset),
    .io_in_0_ready(acqArb_io_in_0_ready),
    .io_in_0_valid(acqArb_io_in_0_valid),
    .io_in_0_bits_addr_block(acqArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(acqArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(acqArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(acqArb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(acqArb_io_in_0_bits_a_type),
    .io_in_0_bits_union(acqArb_io_in_0_bits_union),
    .io_in_0_bits_data(acqArb_io_in_0_bits_data),
    .io_in_1_ready(acqArb_io_in_1_ready),
    .io_in_1_valid(acqArb_io_in_1_valid),
    .io_in_1_bits_addr_block(acqArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(acqArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(acqArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(acqArb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(acqArb_io_in_1_bits_a_type),
    .io_in_1_bits_union(acqArb_io_in_1_bits_union),
    .io_in_1_bits_data(acqArb_io_in_1_bits_data),
    .io_out_ready(acqArb_io_out_ready),
    .io_out_valid(acqArb_io_out_valid),
    .io_out_bits_addr_block(acqArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(acqArb_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(acqArb_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(acqArb_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(acqArb_io_out_bits_a_type),
    .io_out_bits_union(acqArb_io_out_bits_union),
    .io_out_bits_data(acqArb_io_out_bits_data),
    .io_chosen(acqArb_io_chosen)
  );
  ReorderQueue acqRoq (
    .clk(acqRoq_clk),
    .reset(acqRoq_reset),
    .io_enq_ready(acqRoq_io_enq_ready),
    .io_enq_valid(acqRoq_io_enq_valid),
    .io_enq_bits_data(acqRoq_io_enq_bits_data),
    .io_enq_bits_tag(acqRoq_io_enq_bits_tag),
    .io_deq_valid(acqRoq_io_deq_valid),
    .io_deq_tag(acqRoq_io_deq_tag),
    .io_deq_data(acqRoq_io_deq_data),
    .io_deq_matches(acqRoq_io_deq_matches)
  );
  ReorderQueue relRoq (
    .clk(relRoq_clk),
    .reset(relRoq_reset),
    .io_enq_ready(relRoq_io_enq_ready),
    .io_enq_valid(relRoq_io_enq_valid),
    .io_enq_bits_data(relRoq_io_enq_bits_data),
    .io_enq_bits_tag(relRoq_io_enq_bits_tag),
    .io_deq_valid(relRoq_io_deq_valid),
    .io_deq_tag(relRoq_io_deq_tag),
    .io_deq_data(relRoq_io_deq_data),
    .io_deq_matches(relRoq_io_deq_matches)
  );
  assign io_in_acquire_ready = T_1451;
  assign io_in_probe_valid = 1'h0;
  assign io_in_probe_bits_addr_block = GEN_1;
  assign io_in_probe_bits_p_type = GEN_2;
  assign io_in_release_ready = T_1605;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_grant_bits_addr_beat = T_1751_addr_beat;
  assign io_in_grant_bits_client_xact_id = T_1751_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = T_1751_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = T_1751_is_builtin_type;
  assign io_in_grant_bits_g_type = T_1751_g_type;
  assign io_in_grant_bits_data = T_1751_data;
  assign io_in_grant_bits_manager_id = GEN_3;
  assign io_in_finish_ready = 1'h0;
  assign io_out_acquire_valid = acqArb_io_out_valid;
  assign io_out_acquire_bits_addr_block = acqArb_io_out_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = acqArb_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = acqArb_io_out_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = acqArb_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = acqArb_io_out_bits_a_type;
  assign io_out_acquire_bits_union = acqArb_io_out_bits_union;
  assign io_out_acquire_bits_data = acqArb_io_out_bits_data;
  assign io_out_grant_ready = io_in_grant_ready;
  assign acqArb_clk = clk;
  assign acqArb_reset = reset;
  assign acqArb_io_in_0_valid = T_1391;
  assign acqArb_io_in_0_bits_addr_block = T_1423_addr_block;
  assign acqArb_io_in_0_bits_client_xact_id = T_1423_client_xact_id;
  assign acqArb_io_in_0_bits_addr_beat = T_1423_addr_beat;
  assign acqArb_io_in_0_bits_is_builtin_type = T_1423_is_builtin_type;
  assign acqArb_io_in_0_bits_a_type = T_1423_a_type;
  assign acqArb_io_in_0_bits_union = T_1423_union;
  assign acqArb_io_in_0_bits_data = T_1423_data;
  assign acqArb_io_in_1_valid = T_1454;
  assign acqArb_io_in_1_bits_addr_block = T_1577_addr_block;
  assign acqArb_io_in_1_bits_client_xact_id = T_1577_client_xact_id;
  assign acqArb_io_in_1_bits_addr_beat = T_1577_addr_beat;
  assign acqArb_io_in_1_bits_is_builtin_type = T_1577_is_builtin_type;
  assign acqArb_io_in_1_bits_a_type = T_1577_a_type;
  assign acqArb_io_in_1_bits_union = T_1577_union;
  assign acqArb_io_in_1_bits_data = T_1577_data;
  assign acqArb_io_out_ready = io_out_acquire_ready;
  assign acqRoq_clk = clk;
  assign acqRoq_reset = reset;
  assign acqRoq_io_enq_valid = T_1390;
  assign acqRoq_io_enq_bits_data = io_in_acquire_bits_is_builtin_type;
  assign acqRoq_io_enq_bits_tag = io_in_acquire_bits_client_xact_id;
  assign acqRoq_io_deq_valid = T_1625;
  assign acqRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign relRoq_clk = clk;
  assign relRoq_reset = reset;
  assign relRoq_io_enq_valid = T_1453;
  assign relRoq_io_enq_bits_data = io_in_release_bits_voluntary;
  assign relRoq_io_enq_bits_tag = io_in_release_bits_client_xact_id;
  assign relRoq_io_deq_valid = T_1628;
  assign relRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign T_1366_0 = 3'h3;
  assign T_1368 = io_in_acquire_bits_a_type == T_1366_0;
  assign T_1369 = io_in_acquire_bits_is_builtin_type & T_1368;
  assign T_1371 = T_1369 == 1'h0;
  assign T_1373 = io_in_acquire_bits_addr_beat == 3'h0;
  assign acq_roq_enq = T_1371 | T_1373;
  assign T_1375 = io_in_release_bits_r_type == 3'h0;
  assign T_1376 = io_in_release_bits_r_type == 3'h1;
  assign T_1377 = io_in_release_bits_r_type == 3'h2;
  assign T_1378 = T_1375 | T_1376;
  assign T_1379 = T_1378 | T_1377;
  assign T_1382 = T_1379 == 1'h0;
  assign T_1384 = io_in_release_bits_addr_beat == 3'h0;
  assign rel_roq_enq = T_1382 | T_1384;
  assign T_1386 = acq_roq_enq == 1'h0;
  assign acq_roq_ready = T_1386 | acqRoq_io_enq_ready;
  assign T_1388 = rel_roq_enq == 1'h0;
  assign rel_roq_ready = T_1388 | relRoq_io_enq_ready;
  assign T_1389 = io_in_acquire_valid & acqArb_io_in_0_ready;
  assign T_1390 = T_1389 & acq_roq_enq;
  assign T_1391 = io_in_acquire_valid & acq_roq_ready;
  assign T_1394 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_a_type : 3'h1;
  assign T_1423_addr_block = io_in_acquire_bits_addr_block;
  assign T_1423_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign T_1423_addr_beat = io_in_acquire_bits_addr_beat;
  assign T_1423_is_builtin_type = 1'h1;
  assign T_1423_a_type = T_1394;
  assign T_1423_union = io_in_acquire_bits_union;
  assign T_1423_data = io_in_acquire_bits_data;
  assign T_1451 = acq_roq_ready & acqArb_io_in_0_ready;
  assign T_1452 = io_in_release_valid & acqArb_io_in_1_ready;
  assign T_1453 = T_1452 & rel_roq_enq;
  assign T_1454 = io_in_release_valid & rel_roq_ready;
  assign T_1577_addr_block = io_in_release_bits_addr_block;
  assign T_1577_client_xact_id = io_in_release_bits_client_xact_id;
  assign T_1577_addr_beat = io_in_release_bits_addr_beat;
  assign T_1577_is_builtin_type = 1'h1;
  assign T_1577_a_type = 3'h3;
  assign T_1577_union = 11'h1ff;
  assign T_1577_data = io_in_release_bits_data;
  assign T_1605 = rel_roq_ready & acqArb_io_in_1_ready;
  assign T_1606 = io_out_grant_ready & io_out_grant_valid;
  assign T_1614_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_1614_0};
  assign T_1616 = io_out_grant_bits_g_type == GEN_0;
  assign T_1617 = io_out_grant_bits_g_type == 4'h0;
  assign T_1618 = io_out_grant_bits_is_builtin_type ? T_1616 : T_1617;
  assign T_1621 = T_1618 == 1'h0;
  assign T_1623 = io_out_grant_bits_addr_beat == 3'h7;
  assign T_1624 = T_1621 | T_1623;
  assign grant_deq_roq = T_1606 & T_1624;
  assign T_1625 = acqRoq_io_deq_matches & grant_deq_roq;
  assign T_1627 = acqRoq_io_deq_matches == 1'h0;
  assign T_1628 = T_1627 & grant_deq_roq;
  assign T_1630 = grant_deq_roq == 1'h0;
  assign T_1631 = T_1630 | acqRoq_io_deq_matches;
  assign T_1632 = T_1631 | relRoq_io_deq_matches;
  assign T_1633 = T_1632 | reset;
  assign T_1635 = T_1633 == 1'h0;
  assign T_1636 = acqRoq_io_deq_data ? io_out_grant_bits_g_type : 4'h0;
  assign acq_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign acq_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign acq_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign acq_grant_is_builtin_type = acqRoq_io_deq_data;
  assign acq_grant_g_type = T_1636;
  assign acq_grant_data = io_out_grant_bits_data;
  assign T_1691 = io_in_release_valid == 1'h0;
  assign T_1692 = T_1691 | io_in_release_bits_voluntary;
  assign T_1693 = T_1692 | reset;
  assign T_1695 = T_1693 == 1'h0;
  assign rel_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign rel_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign rel_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign rel_grant_is_builtin_type = 1'h1;
  assign rel_grant_g_type = 4'h0;
  assign rel_grant_data = io_out_grant_bits_data;
  assign T_1751_addr_beat = acqRoq_io_deq_matches ? acq_grant_addr_beat : rel_grant_addr_beat;
  assign T_1751_client_xact_id = acqRoq_io_deq_matches ? acq_grant_client_xact_id : rel_grant_client_xact_id;
  assign T_1751_manager_xact_id = acqRoq_io_deq_matches ? acq_grant_manager_xact_id : rel_grant_manager_xact_id;
  assign T_1751_is_builtin_type = acqRoq_io_deq_matches ? acq_grant_is_builtin_type : rel_grant_is_builtin_type;
  assign T_1751_g_type = acqRoq_io_deq_matches ? acq_grant_g_type : rel_grant_g_type;
  assign T_1751_data = acqRoq_io_deq_matches ? acq_grant_data : rel_grant_data;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_4[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_5[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_6[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_4 = {1{$random}};
  GEN_5 = {1{$random}};
  GEN_6 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1635) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink Unwrapper: client_xact_id mismatch\n    at Tilelink.scala:120 assert(!grant_deq_roq || acqRoq.io.deq.matches || relRoq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1635) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1695) begin
          $fwrite(32'h80000002,"Assertion failed: Unwrapper can only process voluntary releases.\n    at Tilelink.scala:134 assert(!io.in.release.valid || io.in.release.bits.isVoluntary(), \"Unwrapper can only process voluntary releases.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1695) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientTileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output  io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_manager_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input   io_inner_finish_bits_manager_xact_id,
  input   io_inner_finish_bits_manager_id,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [1:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id
);
  assign io_inner_acquire_ready = io_outer_acquire_ready;
  assign io_inner_probe_valid = io_outer_probe_valid;
  assign io_inner_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign io_inner_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign io_inner_release_ready = io_outer_release_ready;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_manager_id = io_outer_grant_bits_manager_id;
  assign io_inner_finish_ready = io_outer_finish_ready;
  assign io_outer_acquire_valid = io_inner_acquire_valid;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_probe_ready = io_inner_probe_ready;
  assign io_outer_release_valid = io_inner_release_valid;
  assign io_outer_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign io_outer_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign io_outer_release_bits_r_type = io_inner_release_bits_r_type;
  assign io_outer_release_bits_data = io_inner_release_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_finish_valid = io_inner_finish_valid;
  assign io_outer_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign io_outer_finish_bits_manager_id = io_inner_finish_bits_manager_id;
endmodule
module Queue_10(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [25:0] io_enq_bits_addr_block,
  input   io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input  [10:0] io_enq_bits_union,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [25:0] io_deq_bits_addr_block,
  output  io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [10:0] io_deq_bits_union,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [25:0] ram_addr_block [0:0];
  reg [31:0] GEN_0;
  wire [25:0] ram_addr_block_T_304_data;
  wire  ram_addr_block_T_304_addr;
  wire  ram_addr_block_T_304_en;
  wire [25:0] ram_addr_block_T_269_data;
  wire  ram_addr_block_T_269_addr;
  wire  ram_addr_block_T_269_mask;
  wire  ram_addr_block_T_269_en;
  reg  ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire  ram_client_xact_id_T_304_data;
  wire  ram_client_xact_id_T_304_addr;
  wire  ram_client_xact_id_T_304_en;
  wire  ram_client_xact_id_T_269_data;
  wire  ram_client_xact_id_T_269_addr;
  wire  ram_client_xact_id_T_269_mask;
  wire  ram_client_xact_id_T_269_en;
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_addr_beat_T_304_data;
  wire  ram_addr_beat_T_304_addr;
  wire  ram_addr_beat_T_304_en;
  wire [2:0] ram_addr_beat_T_269_data;
  wire  ram_addr_beat_T_269_addr;
  wire  ram_addr_beat_T_269_mask;
  wire  ram_addr_beat_T_269_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_304_data;
  wire  ram_is_builtin_type_T_304_addr;
  wire  ram_is_builtin_type_T_304_en;
  wire  ram_is_builtin_type_T_269_data;
  wire  ram_is_builtin_type_T_269_addr;
  wire  ram_is_builtin_type_T_269_mask;
  wire  ram_is_builtin_type_T_269_en;
  reg [2:0] ram_a_type [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_304_data;
  wire  ram_a_type_T_304_addr;
  wire  ram_a_type_T_304_en;
  wire [2:0] ram_a_type_T_269_data;
  wire  ram_a_type_T_269_addr;
  wire  ram_a_type_T_269_mask;
  wire  ram_a_type_T_269_en;
  reg [10:0] ram_union [0:0];
  reg [31:0] GEN_5;
  wire [10:0] ram_union_T_304_data;
  wire  ram_union_T_304_addr;
  wire  ram_union_T_304_en;
  wire [10:0] ram_union_T_269_data;
  wire  ram_union_T_269_addr;
  wire  ram_union_T_269_mask;
  wire  ram_union_T_269_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_6;
  wire [63:0] ram_data_T_304_data;
  wire  ram_data_T_304_addr;
  wire  ram_data_T_304_en;
  wire [63:0] ram_data_T_269_data;
  wire  ram_data_T_269_addr;
  wire  ram_data_T_269_mask;
  wire  ram_data_T_269_en;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  T_266;
  wire  T_267;
  wire  do_enq;
  wire  T_268;
  wire  do_deq;
  wire  T_299;
  wire  GEN_17;
  wire  T_301;
  wire [1:0] T_332;
  wire  ptr_diff;
  wire [1:0] T_334;
  assign io_enq_ready = T_266;
  assign io_deq_valid = T_301;
  assign io_deq_bits_addr_block = ram_addr_block_T_304_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_304_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_304_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_304_data;
  assign io_deq_bits_a_type = ram_a_type_T_304_data;
  assign io_deq_bits_union = ram_union_T_304_data;
  assign io_deq_bits_data = ram_data_T_304_data;
  assign io_count = T_334[0];
  assign ram_addr_block_T_304_addr = 1'h0;
  assign ram_addr_block_T_304_en = 1'h1;
  assign ram_addr_block_T_304_data = ram_addr_block[ram_addr_block_T_304_addr];
  assign ram_addr_block_T_269_data = io_enq_bits_addr_block;
  assign ram_addr_block_T_269_addr = 1'h0;
  assign ram_addr_block_T_269_mask = do_enq;
  assign ram_addr_block_T_269_en = do_enq;
  assign ram_client_xact_id_T_304_addr = 1'h0;
  assign ram_client_xact_id_T_304_en = 1'h1;
  assign ram_client_xact_id_T_304_data = ram_client_xact_id[ram_client_xact_id_T_304_addr];
  assign ram_client_xact_id_T_269_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_269_addr = 1'h0;
  assign ram_client_xact_id_T_269_mask = do_enq;
  assign ram_client_xact_id_T_269_en = do_enq;
  assign ram_addr_beat_T_304_addr = 1'h0;
  assign ram_addr_beat_T_304_en = 1'h1;
  assign ram_addr_beat_T_304_data = ram_addr_beat[ram_addr_beat_T_304_addr];
  assign ram_addr_beat_T_269_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_269_addr = 1'h0;
  assign ram_addr_beat_T_269_mask = do_enq;
  assign ram_addr_beat_T_269_en = do_enq;
  assign ram_is_builtin_type_T_304_addr = 1'h0;
  assign ram_is_builtin_type_T_304_en = 1'h1;
  assign ram_is_builtin_type_T_304_data = ram_is_builtin_type[ram_is_builtin_type_T_304_addr];
  assign ram_is_builtin_type_T_269_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_269_addr = 1'h0;
  assign ram_is_builtin_type_T_269_mask = do_enq;
  assign ram_is_builtin_type_T_269_en = do_enq;
  assign ram_a_type_T_304_addr = 1'h0;
  assign ram_a_type_T_304_en = 1'h1;
  assign ram_a_type_T_304_data = ram_a_type[ram_a_type_T_304_addr];
  assign ram_a_type_T_269_data = io_enq_bits_a_type;
  assign ram_a_type_T_269_addr = 1'h0;
  assign ram_a_type_T_269_mask = do_enq;
  assign ram_a_type_T_269_en = do_enq;
  assign ram_union_T_304_addr = 1'h0;
  assign ram_union_T_304_en = 1'h1;
  assign ram_union_T_304_data = ram_union[ram_union_T_304_addr];
  assign ram_union_T_269_data = io_enq_bits_union;
  assign ram_union_T_269_addr = 1'h0;
  assign ram_union_T_269_mask = do_enq;
  assign ram_union_T_269_en = do_enq;
  assign ram_data_T_304_addr = 1'h0;
  assign ram_data_T_304_en = 1'h1;
  assign ram_data_T_304_data = ram_data[ram_data_T_304_addr];
  assign ram_data_T_269_data = io_enq_bits_data;
  assign ram_data_T_269_addr = 1'h0;
  assign ram_data_T_269_mask = do_enq;
  assign ram_data_T_269_en = do_enq;
  assign T_266 = maybe_full == 1'h0;
  assign T_267 = io_enq_ready & io_enq_valid;
  assign do_enq = T_267;
  assign T_268 = io_deq_ready & io_deq_valid;
  assign do_deq = T_268;
  assign T_299 = do_enq != do_deq;
  assign GEN_17 = T_299 ? do_enq : maybe_full;
  assign T_301 = T_266 == 1'h0;
  assign T_332 = 1'h0 - 1'h0;
  assign ptr_diff = T_332[0:0];
  assign T_334 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_block[initvar] = GEN_0[25:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[0:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_union[initvar] = GEN_5[10:0];
  `endif
  GEN_6 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_6[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_block_T_269_en & ram_addr_block_T_269_mask) begin
      ram_addr_block[ram_addr_block_T_269_addr] <= ram_addr_block_T_269_data;
    end
    if(ram_client_xact_id_T_269_en & ram_client_xact_id_T_269_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_269_addr] <= ram_client_xact_id_T_269_data;
    end
    if(ram_addr_beat_T_269_en & ram_addr_beat_T_269_mask) begin
      ram_addr_beat[ram_addr_beat_T_269_addr] <= ram_addr_beat_T_269_data;
    end
    if(ram_is_builtin_type_T_269_en & ram_is_builtin_type_T_269_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_269_addr] <= ram_is_builtin_type_T_269_data;
    end
    if(ram_a_type_T_269_en & ram_a_type_T_269_mask) begin
      ram_a_type[ram_a_type_T_269_addr] <= ram_a_type_T_269_data;
    end
    if(ram_union_T_269_en & ram_union_T_269_mask) begin
      ram_union[ram_union_T_269_addr] <= ram_union_T_269_data;
    end
    if(ram_data_T_269_en & ram_data_T_269_mask) begin
      ram_data[ram_data_T_269_addr] <= ram_data_T_269_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_299) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_11(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_client_xact_id,
  input  [1:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_is_builtin_type,
  input  [3:0] io_enq_bits_g_type,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_client_xact_id,
  output [1:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_is_builtin_type,
  output [3:0] io_deq_bits_g_type,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_0;
  wire [2:0] ram_addr_beat_T_294_data;
  wire  ram_addr_beat_T_294_addr;
  wire  ram_addr_beat_T_294_en;
  wire [2:0] ram_addr_beat_T_260_data;
  wire  ram_addr_beat_T_260_addr;
  wire  ram_addr_beat_T_260_mask;
  wire  ram_addr_beat_T_260_en;
  reg  ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire  ram_client_xact_id_T_294_data;
  wire  ram_client_xact_id_T_294_addr;
  wire  ram_client_xact_id_T_294_en;
  wire  ram_client_xact_id_T_260_data;
  wire  ram_client_xact_id_T_260_addr;
  wire  ram_client_xact_id_T_260_mask;
  wire  ram_client_xact_id_T_260_en;
  reg [1:0] ram_manager_xact_id [0:0];
  reg [31:0] GEN_2;
  wire [1:0] ram_manager_xact_id_T_294_data;
  wire  ram_manager_xact_id_T_294_addr;
  wire  ram_manager_xact_id_T_294_en;
  wire [1:0] ram_manager_xact_id_T_260_data;
  wire  ram_manager_xact_id_T_260_addr;
  wire  ram_manager_xact_id_T_260_mask;
  wire  ram_manager_xact_id_T_260_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_294_data;
  wire  ram_is_builtin_type_T_294_addr;
  wire  ram_is_builtin_type_T_294_en;
  wire  ram_is_builtin_type_T_260_data;
  wire  ram_is_builtin_type_T_260_addr;
  wire  ram_is_builtin_type_T_260_mask;
  wire  ram_is_builtin_type_T_260_en;
  reg [3:0] ram_g_type [0:0];
  reg [31:0] GEN_4;
  wire [3:0] ram_g_type_T_294_data;
  wire  ram_g_type_T_294_addr;
  wire  ram_g_type_T_294_en;
  wire [3:0] ram_g_type_T_260_data;
  wire  ram_g_type_T_260_addr;
  wire  ram_g_type_T_260_mask;
  wire  ram_g_type_T_260_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_5;
  wire [63:0] ram_data_T_294_data;
  wire  ram_data_T_294_addr;
  wire  ram_data_T_294_en;
  wire [63:0] ram_data_T_260_data;
  wire  ram_data_T_260_addr;
  wire  ram_data_T_260_mask;
  wire  ram_data_T_260_en;
  reg  maybe_full;
  reg [31:0] GEN_6;
  wire  T_257;
  wire  T_258;
  wire  do_enq;
  wire  T_259;
  wire  do_deq;
  wire  T_289;
  wire  GEN_15;
  wire  T_291;
  wire [1:0] T_321;
  wire  ptr_diff;
  wire [1:0] T_323;
  assign io_enq_ready = T_257;
  assign io_deq_valid = T_291;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_294_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_294_data;
  assign io_deq_bits_manager_xact_id = ram_manager_xact_id_T_294_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_294_data;
  assign io_deq_bits_g_type = ram_g_type_T_294_data;
  assign io_deq_bits_data = ram_data_T_294_data;
  assign io_count = T_323[0];
  assign ram_addr_beat_T_294_addr = 1'h0;
  assign ram_addr_beat_T_294_en = 1'h1;
  assign ram_addr_beat_T_294_data = ram_addr_beat[ram_addr_beat_T_294_addr];
  assign ram_addr_beat_T_260_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_260_addr = 1'h0;
  assign ram_addr_beat_T_260_mask = do_enq;
  assign ram_addr_beat_T_260_en = do_enq;
  assign ram_client_xact_id_T_294_addr = 1'h0;
  assign ram_client_xact_id_T_294_en = 1'h1;
  assign ram_client_xact_id_T_294_data = ram_client_xact_id[ram_client_xact_id_T_294_addr];
  assign ram_client_xact_id_T_260_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_260_addr = 1'h0;
  assign ram_client_xact_id_T_260_mask = do_enq;
  assign ram_client_xact_id_T_260_en = do_enq;
  assign ram_manager_xact_id_T_294_addr = 1'h0;
  assign ram_manager_xact_id_T_294_en = 1'h1;
  assign ram_manager_xact_id_T_294_data = ram_manager_xact_id[ram_manager_xact_id_T_294_addr];
  assign ram_manager_xact_id_T_260_data = io_enq_bits_manager_xact_id;
  assign ram_manager_xact_id_T_260_addr = 1'h0;
  assign ram_manager_xact_id_T_260_mask = do_enq;
  assign ram_manager_xact_id_T_260_en = do_enq;
  assign ram_is_builtin_type_T_294_addr = 1'h0;
  assign ram_is_builtin_type_T_294_en = 1'h1;
  assign ram_is_builtin_type_T_294_data = ram_is_builtin_type[ram_is_builtin_type_T_294_addr];
  assign ram_is_builtin_type_T_260_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_260_addr = 1'h0;
  assign ram_is_builtin_type_T_260_mask = do_enq;
  assign ram_is_builtin_type_T_260_en = do_enq;
  assign ram_g_type_T_294_addr = 1'h0;
  assign ram_g_type_T_294_en = 1'h1;
  assign ram_g_type_T_294_data = ram_g_type[ram_g_type_T_294_addr];
  assign ram_g_type_T_260_data = io_enq_bits_g_type;
  assign ram_g_type_T_260_addr = 1'h0;
  assign ram_g_type_T_260_mask = do_enq;
  assign ram_g_type_T_260_en = do_enq;
  assign ram_data_T_294_addr = 1'h0;
  assign ram_data_T_294_en = 1'h1;
  assign ram_data_T_294_data = ram_data[ram_data_T_294_addr];
  assign ram_data_T_260_data = io_enq_bits_data;
  assign ram_data_T_260_addr = 1'h0;
  assign ram_data_T_260_mask = do_enq;
  assign ram_data_T_260_en = do_enq;
  assign T_257 = maybe_full == 1'h0;
  assign T_258 = io_enq_ready & io_enq_valid;
  assign do_enq = T_258;
  assign T_259 = io_deq_ready & io_deq_valid;
  assign do_deq = T_259;
  assign T_289 = do_enq != do_deq;
  assign GEN_15 = T_289 ? do_enq : maybe_full;
  assign T_291 = T_257 == 1'h0;
  assign T_321 = 1'h0 - 1'h0;
  assign ptr_diff = T_321[0:0];
  assign T_323 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_0[2:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[0:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_manager_xact_id[initvar] = GEN_2[1:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_g_type[initvar] = GEN_4[3:0];
  `endif
  GEN_5 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_5[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  maybe_full = GEN_6[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_beat_T_260_en & ram_addr_beat_T_260_mask) begin
      ram_addr_beat[ram_addr_beat_T_260_addr] <= ram_addr_beat_T_260_data;
    end
    if(ram_client_xact_id_T_260_en & ram_client_xact_id_T_260_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_260_addr] <= ram_client_xact_id_T_260_data;
    end
    if(ram_manager_xact_id_T_260_en & ram_manager_xact_id_T_260_mask) begin
      ram_manager_xact_id[ram_manager_xact_id_T_260_addr] <= ram_manager_xact_id_T_260_data;
    end
    if(ram_is_builtin_type_T_260_en & ram_is_builtin_type_T_260_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_260_addr] <= ram_is_builtin_type_T_260_data;
    end
    if(ram_g_type_T_260_en & ram_g_type_T_260_mask) begin
      ram_g_type[ram_g_type_T_260_addr] <= ram_g_type_T_260_data;
    end
    if(ram_data_T_260_en & ram_data_T_260_mask) begin
      ram_data[ram_data_T_260_addr] <= ram_data_T_260_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_289) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module ClientUncachedTileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input   io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output  io_inner_grant_bits_client_xact_id,
  output [1:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output  io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input   io_outer_grant_bits_client_xact_id,
  input  [1:0] io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data
);
  wire  Queue_10_1_clk;
  wire  Queue_10_1_reset;
  wire  Queue_10_1_io_enq_ready;
  wire  Queue_10_1_io_enq_valid;
  wire [25:0] Queue_10_1_io_enq_bits_addr_block;
  wire  Queue_10_1_io_enq_bits_client_xact_id;
  wire [2:0] Queue_10_1_io_enq_bits_addr_beat;
  wire  Queue_10_1_io_enq_bits_is_builtin_type;
  wire [2:0] Queue_10_1_io_enq_bits_a_type;
  wire [10:0] Queue_10_1_io_enq_bits_union;
  wire [63:0] Queue_10_1_io_enq_bits_data;
  wire  Queue_10_1_io_deq_ready;
  wire  Queue_10_1_io_deq_valid;
  wire [25:0] Queue_10_1_io_deq_bits_addr_block;
  wire  Queue_10_1_io_deq_bits_client_xact_id;
  wire [2:0] Queue_10_1_io_deq_bits_addr_beat;
  wire  Queue_10_1_io_deq_bits_is_builtin_type;
  wire [2:0] Queue_10_1_io_deq_bits_a_type;
  wire [10:0] Queue_10_1_io_deq_bits_union;
  wire [63:0] Queue_10_1_io_deq_bits_data;
  wire  Queue_10_1_io_count;
  wire  Queue_11_1_clk;
  wire  Queue_11_1_reset;
  wire  Queue_11_1_io_enq_ready;
  wire  Queue_11_1_io_enq_valid;
  wire [2:0] Queue_11_1_io_enq_bits_addr_beat;
  wire  Queue_11_1_io_enq_bits_client_xact_id;
  wire [1:0] Queue_11_1_io_enq_bits_manager_xact_id;
  wire  Queue_11_1_io_enq_bits_is_builtin_type;
  wire [3:0] Queue_11_1_io_enq_bits_g_type;
  wire [63:0] Queue_11_1_io_enq_bits_data;
  wire  Queue_11_1_io_deq_ready;
  wire  Queue_11_1_io_deq_valid;
  wire [2:0] Queue_11_1_io_deq_bits_addr_beat;
  wire  Queue_11_1_io_deq_bits_client_xact_id;
  wire [1:0] Queue_11_1_io_deq_bits_manager_xact_id;
  wire  Queue_11_1_io_deq_bits_is_builtin_type;
  wire [3:0] Queue_11_1_io_deq_bits_g_type;
  wire [63:0] Queue_11_1_io_deq_bits_data;
  wire  Queue_11_1_io_count;
  Queue_10 Queue_10_1 (
    .clk(Queue_10_1_clk),
    .reset(Queue_10_1_reset),
    .io_enq_ready(Queue_10_1_io_enq_ready),
    .io_enq_valid(Queue_10_1_io_enq_valid),
    .io_enq_bits_addr_block(Queue_10_1_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(Queue_10_1_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(Queue_10_1_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(Queue_10_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(Queue_10_1_io_enq_bits_a_type),
    .io_enq_bits_union(Queue_10_1_io_enq_bits_union),
    .io_enq_bits_data(Queue_10_1_io_enq_bits_data),
    .io_deq_ready(Queue_10_1_io_deq_ready),
    .io_deq_valid(Queue_10_1_io_deq_valid),
    .io_deq_bits_addr_block(Queue_10_1_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(Queue_10_1_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(Queue_10_1_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(Queue_10_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(Queue_10_1_io_deq_bits_a_type),
    .io_deq_bits_union(Queue_10_1_io_deq_bits_union),
    .io_deq_bits_data(Queue_10_1_io_deq_bits_data),
    .io_count(Queue_10_1_io_count)
  );
  Queue_11 Queue_11_1 (
    .clk(Queue_11_1_clk),
    .reset(Queue_11_1_reset),
    .io_enq_ready(Queue_11_1_io_enq_ready),
    .io_enq_valid(Queue_11_1_io_enq_valid),
    .io_enq_bits_addr_beat(Queue_11_1_io_enq_bits_addr_beat),
    .io_enq_bits_client_xact_id(Queue_11_1_io_enq_bits_client_xact_id),
    .io_enq_bits_manager_xact_id(Queue_11_1_io_enq_bits_manager_xact_id),
    .io_enq_bits_is_builtin_type(Queue_11_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_g_type(Queue_11_1_io_enq_bits_g_type),
    .io_enq_bits_data(Queue_11_1_io_enq_bits_data),
    .io_deq_ready(Queue_11_1_io_deq_ready),
    .io_deq_valid(Queue_11_1_io_deq_valid),
    .io_deq_bits_addr_beat(Queue_11_1_io_deq_bits_addr_beat),
    .io_deq_bits_client_xact_id(Queue_11_1_io_deq_bits_client_xact_id),
    .io_deq_bits_manager_xact_id(Queue_11_1_io_deq_bits_manager_xact_id),
    .io_deq_bits_is_builtin_type(Queue_11_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_g_type(Queue_11_1_io_deq_bits_g_type),
    .io_deq_bits_data(Queue_11_1_io_deq_bits_data),
    .io_count(Queue_11_1_io_count)
  );
  assign io_inner_acquire_ready = Queue_10_1_io_enq_ready;
  assign io_inner_grant_valid = Queue_11_1_io_deq_valid;
  assign io_inner_grant_bits_addr_beat = Queue_11_1_io_deq_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = Queue_11_1_io_deq_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = Queue_11_1_io_deq_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = Queue_11_1_io_deq_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = Queue_11_1_io_deq_bits_g_type;
  assign io_inner_grant_bits_data = Queue_11_1_io_deq_bits_data;
  assign io_outer_acquire_valid = Queue_10_1_io_deq_valid;
  assign io_outer_acquire_bits_addr_block = Queue_10_1_io_deq_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = Queue_10_1_io_deq_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = Queue_10_1_io_deq_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = Queue_10_1_io_deq_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = Queue_10_1_io_deq_bits_a_type;
  assign io_outer_acquire_bits_union = Queue_10_1_io_deq_bits_union;
  assign io_outer_acquire_bits_data = Queue_10_1_io_deq_bits_data;
  assign io_outer_grant_ready = Queue_11_1_io_enq_ready;
  assign Queue_10_1_clk = clk;
  assign Queue_10_1_reset = reset;
  assign Queue_10_1_io_enq_valid = io_inner_acquire_valid;
  assign Queue_10_1_io_enq_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign Queue_10_1_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign Queue_10_1_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign Queue_10_1_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign Queue_10_1_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign Queue_10_1_io_enq_bits_union = io_inner_acquire_bits_union;
  assign Queue_10_1_io_enq_bits_data = io_inner_acquire_bits_data;
  assign Queue_10_1_io_deq_ready = io_outer_acquire_ready;
  assign Queue_11_1_clk = clk;
  assign Queue_11_1_reset = reset;
  assign Queue_11_1_io_enq_valid = io_outer_grant_valid;
  assign Queue_11_1_io_enq_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign Queue_11_1_io_enq_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign Queue_11_1_io_enq_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign Queue_11_1_io_enq_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign Queue_11_1_io_enq_bits_g_type = io_outer_grant_bits_g_type;
  assign Queue_11_1_io_enq_bits_data = io_outer_grant_bits_data;
  assign Queue_11_1_io_deq_ready = io_inner_grant_ready;
endmodule
module LockingRRArbiter_10(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire  GEN_0_bits_manager_xact_id;
  wire  GEN_0_bits_is_builtin_type;
  wire [3:0] GEN_0_bits_g_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire  GEN_1_bits_manager_xact_id;
  wire  GEN_1_bits_is_builtin_type;
  wire [3:0] GEN_1_bits_g_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire  GEN_2_bits_manager_xact_id;
  wire  GEN_2_bits_is_builtin_type;
  wire [3:0] GEN_2_bits_g_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire  GEN_3_bits_manager_xact_id;
  wire  GEN_3_bits_is_builtin_type;
  wire [3:0] GEN_3_bits_g_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire  GEN_4_bits_manager_xact_id;
  wire  GEN_4_bits_is_builtin_type;
  wire [3:0] GEN_4_bits_g_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire  GEN_5_bits_manager_xact_id;
  wire  GEN_5_bits_is_builtin_type;
  wire [3:0] GEN_5_bits_g_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire  GEN_6_bits_manager_xact_id;
  wire  GEN_6_bits_is_builtin_type;
  wire [3:0] GEN_6_bits_g_type;
  wire [63:0] GEN_6_bits_data;
  reg [2:0] T_518;
  reg [31:0] GEN_1;
  reg  T_520;
  reg [31:0] GEN_2;
  wire  T_522;
  wire [2:0] T_530_0;
  wire [3:0] GEN_0;
  wire  T_532;
  wire  T_533;
  wire  T_534;
  wire  T_536;
  wire  T_537;
  wire [3:0] T_541;
  wire [2:0] T_542;
  wire  GEN_7;
  wire [2:0] GEN_8;
  wire  GEN_9;
  reg  lastGrant;
  reg [31:0] GEN_3;
  wire  GEN_10;
  wire  T_551;
  wire  T_552;
  wire  T_553;
  assign io_in_0_ready = T_553;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = GEN_3_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_g_type = GEN_5_bits_g_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_chosen = GEN_9;
  assign choice = 1'h0;
  assign GEN_0_ready = io_in_0_ready;
  assign GEN_0_valid = io_in_0_valid;
  assign GEN_0_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_0_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_0_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_0_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_0_bits_g_type = io_in_0_bits_g_type;
  assign GEN_0_bits_data = io_in_0_bits_data;
  assign GEN_1_ready = io_in_0_ready;
  assign GEN_1_valid = io_in_0_valid;
  assign GEN_1_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_1_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_1_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_1_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_1_bits_g_type = io_in_0_bits_g_type;
  assign GEN_1_bits_data = io_in_0_bits_data;
  assign GEN_2_ready = io_in_0_ready;
  assign GEN_2_valid = io_in_0_valid;
  assign GEN_2_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_2_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_2_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_2_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_2_bits_g_type = io_in_0_bits_g_type;
  assign GEN_2_bits_data = io_in_0_bits_data;
  assign GEN_3_ready = io_in_0_ready;
  assign GEN_3_valid = io_in_0_valid;
  assign GEN_3_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_3_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_3_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_3_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_3_bits_g_type = io_in_0_bits_g_type;
  assign GEN_3_bits_data = io_in_0_bits_data;
  assign GEN_4_ready = io_in_0_ready;
  assign GEN_4_valid = io_in_0_valid;
  assign GEN_4_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_4_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_4_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_4_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_4_bits_g_type = io_in_0_bits_g_type;
  assign GEN_4_bits_data = io_in_0_bits_data;
  assign GEN_5_ready = io_in_0_ready;
  assign GEN_5_valid = io_in_0_valid;
  assign GEN_5_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_5_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_5_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_5_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_5_bits_g_type = io_in_0_bits_g_type;
  assign GEN_5_bits_data = io_in_0_bits_data;
  assign GEN_6_ready = io_in_0_ready;
  assign GEN_6_valid = io_in_0_valid;
  assign GEN_6_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_6_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_6_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_6_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_6_bits_g_type = io_in_0_bits_g_type;
  assign GEN_6_bits_data = io_in_0_bits_data;
  assign T_522 = T_518 != 3'h0;
  assign T_530_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_530_0};
  assign T_532 = io_out_bits_g_type == GEN_0;
  assign T_533 = io_out_bits_g_type == 4'h0;
  assign T_534 = io_out_bits_is_builtin_type ? T_532 : T_533;
  assign T_536 = io_out_ready & io_out_valid;
  assign T_537 = T_536 & T_534;
  assign T_541 = T_518 + 3'h1;
  assign T_542 = T_541[2:0];
  assign GEN_7 = T_537 ? io_chosen : T_520;
  assign GEN_8 = T_537 ? T_542 : T_518;
  assign GEN_9 = T_522 ? T_520 : choice;
  assign GEN_10 = T_536 ? io_chosen : lastGrant;
  assign T_551 = T_520 == 1'h0;
  assign T_552 = T_522 ? T_551 : 1'h1;
  assign T_553 = T_552 & io_out_ready;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_518 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_520 = GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  lastGrant = GEN_3[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_518 <= 3'h0;
    end else begin
      if(T_537) begin
        T_518 <= T_542;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_537) begin
        T_520 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_536) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIORouter(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [10:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data
);
  wire [2:0] T_1246_0;
  wire [2:0] T_1246_1;
  wire  T_1248;
  wire  T_1249;
  wire  T_1250;
  wire  T_1251;
  wire [2:0] T_1252;
  wire [2:0] T_1254;
  wire [28:0] T_1255;
  wire [31:0] T_1256;
  wire  T_1260;
  wire  T_1263;
  wire  T_1265;
  wire  T_1266;
  wire  T_1268;
  wire  T_1270;
  wire  T_1271;
  wire  T_1273;
  wire  T_1275;
  wire  T_1276;
  wire  T_1277;
  wire  T_1278;
  wire  acq_route;
  wire  T_1281;
  wire  GEN_0;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_chosen;
  wire  T_1306;
  wire  T_1309;
  wire  T_1310;
  wire  T_1312;
  LockingRRArbiter_10 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_0;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_1281;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign T_1246_0 = 3'h0;
  assign T_1246_1 = 3'h4;
  assign T_1248 = io_in_acquire_bits_a_type == T_1246_0;
  assign T_1249 = io_in_acquire_bits_a_type == T_1246_1;
  assign T_1250 = T_1248 | T_1249;
  assign T_1251 = io_in_acquire_bits_is_builtin_type & T_1250;
  assign T_1252 = io_in_acquire_bits_union[10:8];
  assign T_1254 = T_1251 ? T_1252 : 3'h0;
  assign T_1255 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_1256 = {T_1255,T_1254};
  assign T_1260 = T_1256 < 32'h1000;
  assign T_1263 = 32'h1000 <= T_1256;
  assign T_1265 = T_1256 < 32'h2000;
  assign T_1266 = T_1263 & T_1265;
  assign T_1268 = 32'h40000000 <= T_1256;
  assign T_1270 = T_1256 < 32'h44000000;
  assign T_1271 = T_1268 & T_1270;
  assign T_1273 = 32'h44000000 <= T_1256;
  assign T_1275 = T_1256 < 32'h48000000;
  assign T_1276 = T_1273 & T_1275;
  assign T_1277 = T_1260 | T_1266;
  assign T_1278 = T_1277 | T_1271;
  assign acq_route = T_1278 | T_1276;
  assign T_1281 = io_in_acquire_valid & acq_route;
  assign GEN_0 = acq_route ? io_out_0_acquire_ready : 1'h0;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_1306 = io_in_acquire_valid == 1'h0;
  assign T_1309 = T_1306 | acq_route;
  assign T_1310 = T_1309 | reset;
  assign T_1312 = T_1310 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1312) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at Interconnect.scala:219 assert(!io.in.acquire.valid || acq_route.orR, \"No valid route\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_1_clk;
  wire  ClientUncachedTileLinkIORouter_1_reset;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data;
  ClientUncachedTileLinkIORouter ClientUncachedTileLinkIORouter_1 (
    .clk(ClientUncachedTileLinkIORouter_1_clk),
    .reset(ClientUncachedTileLinkIORouter_1_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_1_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_1_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_1_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_clk = clk;
  assign ClientUncachedTileLinkIORouter_1_reset = reset;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_1_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
endmodule
module LockingRRArbiter_11(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [1:0] io_in_2_bits_client_xact_id,
  input   io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_is_builtin_type,
  input  [3:0] io_in_2_bits_g_type,
  input  [63:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [1:0] io_in_3_bits_client_xact_id,
  input   io_in_3_bits_manager_xact_id,
  input   io_in_3_bits_is_builtin_type,
  input  [3:0] io_in_3_bits_g_type,
  input  [63:0] io_in_3_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire  GEN_0_bits_manager_xact_id;
  wire  GEN_0_bits_is_builtin_type;
  wire [3:0] GEN_0_bits_g_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [1:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [3:0] GEN_13;
  wire [63:0] GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [1:0] GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [3:0] GEN_21;
  wire [63:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [2:0] GEN_25;
  wire [1:0] GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire [3:0] GEN_29;
  wire [63:0] GEN_30;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire  GEN_1_bits_manager_xact_id;
  wire  GEN_1_bits_is_builtin_type;
  wire [3:0] GEN_1_bits_g_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire  GEN_2_bits_manager_xact_id;
  wire  GEN_2_bits_is_builtin_type;
  wire [3:0] GEN_2_bits_g_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire  GEN_3_bits_manager_xact_id;
  wire  GEN_3_bits_is_builtin_type;
  wire [3:0] GEN_3_bits_g_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire  GEN_4_bits_manager_xact_id;
  wire  GEN_4_bits_is_builtin_type;
  wire [3:0] GEN_4_bits_g_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire  GEN_5_bits_manager_xact_id;
  wire  GEN_5_bits_is_builtin_type;
  wire [3:0] GEN_5_bits_g_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire  GEN_6_bits_manager_xact_id;
  wire  GEN_6_bits_is_builtin_type;
  wire [3:0] GEN_6_bits_g_type;
  wire [63:0] GEN_6_bits_data;
  reg [2:0] T_794;
  reg [31:0] GEN_1;
  reg [1:0] T_796;
  reg [31:0] GEN_2;
  wire  T_798;
  wire [2:0] T_806_0;
  wire [3:0] GEN_0;
  wire  T_808;
  wire  T_809;
  wire  T_810;
  wire  T_812;
  wire  T_813;
  wire [3:0] T_817;
  wire [2:0] T_818;
  wire [1:0] GEN_175;
  wire [2:0] GEN_176;
  wire [1:0] GEN_177;
  reg [1:0] lastGrant;
  reg [31:0] GEN_3;
  wire [1:0] GEN_178;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_826;
  wire  T_827;
  wire  T_828;
  wire  T_829;
  wire  T_830;
  wire  T_834;
  wire  T_836;
  wire  T_838;
  wire  T_840;
  wire  T_842;
  wire  T_844;
  wire  T_848;
  wire  T_849;
  wire  T_850;
  wire  T_851;
  wire  T_852;
  wire  T_854;
  wire  T_855;
  wire  T_856;
  wire  T_858;
  wire  T_859;
  wire  T_860;
  wire  T_862;
  wire  T_863;
  wire  T_864;
  wire  T_866;
  wire  T_867;
  wire  T_868;
  wire [1:0] GEN_179;
  wire [1:0] GEN_180;
  wire [1:0] GEN_181;
  wire [1:0] GEN_182;
  wire [1:0] GEN_183;
  wire [1:0] GEN_184;
  assign io_in_0_ready = T_856;
  assign io_in_1_ready = T_860;
  assign io_in_2_ready = T_864;
  assign io_in_3_ready = T_868;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = GEN_3_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_g_type = GEN_5_bits_g_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_chosen = GEN_177;
  assign choice = GEN_184;
  assign GEN_0_ready = GEN_23;
  assign GEN_0_valid = GEN_24;
  assign GEN_0_bits_addr_beat = GEN_25;
  assign GEN_0_bits_client_xact_id = GEN_26;
  assign GEN_0_bits_manager_xact_id = GEN_27;
  assign GEN_0_bits_is_builtin_type = GEN_28;
  assign GEN_0_bits_g_type = GEN_29;
  assign GEN_0_bits_data = GEN_30;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_15 = 2'h2 == io_chosen ? io_in_2_ready : GEN_7;
  assign GEN_16 = 2'h2 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_9;
  assign GEN_18 = 2'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_10;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_manager_xact_id : GEN_11;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_12;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_g_type : GEN_13;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_data : GEN_14;
  assign GEN_23 = 2'h3 == io_chosen ? io_in_3_ready : GEN_15;
  assign GEN_24 = 2'h3 == io_chosen ? io_in_3_valid : GEN_16;
  assign GEN_25 = 2'h3 == io_chosen ? io_in_3_bits_addr_beat : GEN_17;
  assign GEN_26 = 2'h3 == io_chosen ? io_in_3_bits_client_xact_id : GEN_18;
  assign GEN_27 = 2'h3 == io_chosen ? io_in_3_bits_manager_xact_id : GEN_19;
  assign GEN_28 = 2'h3 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_20;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_bits_g_type : GEN_21;
  assign GEN_30 = 2'h3 == io_chosen ? io_in_3_bits_data : GEN_22;
  assign GEN_1_ready = GEN_23;
  assign GEN_1_valid = GEN_24;
  assign GEN_1_bits_addr_beat = GEN_25;
  assign GEN_1_bits_client_xact_id = GEN_26;
  assign GEN_1_bits_manager_xact_id = GEN_27;
  assign GEN_1_bits_is_builtin_type = GEN_28;
  assign GEN_1_bits_g_type = GEN_29;
  assign GEN_1_bits_data = GEN_30;
  assign GEN_2_ready = GEN_23;
  assign GEN_2_valid = GEN_24;
  assign GEN_2_bits_addr_beat = GEN_25;
  assign GEN_2_bits_client_xact_id = GEN_26;
  assign GEN_2_bits_manager_xact_id = GEN_27;
  assign GEN_2_bits_is_builtin_type = GEN_28;
  assign GEN_2_bits_g_type = GEN_29;
  assign GEN_2_bits_data = GEN_30;
  assign GEN_3_ready = GEN_23;
  assign GEN_3_valid = GEN_24;
  assign GEN_3_bits_addr_beat = GEN_25;
  assign GEN_3_bits_client_xact_id = GEN_26;
  assign GEN_3_bits_manager_xact_id = GEN_27;
  assign GEN_3_bits_is_builtin_type = GEN_28;
  assign GEN_3_bits_g_type = GEN_29;
  assign GEN_3_bits_data = GEN_30;
  assign GEN_4_ready = GEN_23;
  assign GEN_4_valid = GEN_24;
  assign GEN_4_bits_addr_beat = GEN_25;
  assign GEN_4_bits_client_xact_id = GEN_26;
  assign GEN_4_bits_manager_xact_id = GEN_27;
  assign GEN_4_bits_is_builtin_type = GEN_28;
  assign GEN_4_bits_g_type = GEN_29;
  assign GEN_4_bits_data = GEN_30;
  assign GEN_5_ready = GEN_23;
  assign GEN_5_valid = GEN_24;
  assign GEN_5_bits_addr_beat = GEN_25;
  assign GEN_5_bits_client_xact_id = GEN_26;
  assign GEN_5_bits_manager_xact_id = GEN_27;
  assign GEN_5_bits_is_builtin_type = GEN_28;
  assign GEN_5_bits_g_type = GEN_29;
  assign GEN_5_bits_data = GEN_30;
  assign GEN_6_ready = GEN_23;
  assign GEN_6_valid = GEN_24;
  assign GEN_6_bits_addr_beat = GEN_25;
  assign GEN_6_bits_client_xact_id = GEN_26;
  assign GEN_6_bits_manager_xact_id = GEN_27;
  assign GEN_6_bits_is_builtin_type = GEN_28;
  assign GEN_6_bits_g_type = GEN_29;
  assign GEN_6_bits_data = GEN_30;
  assign T_798 = T_794 != 3'h0;
  assign T_806_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_806_0};
  assign T_808 = io_out_bits_g_type == GEN_0;
  assign T_809 = io_out_bits_g_type == 4'h0;
  assign T_810 = io_out_bits_is_builtin_type ? T_808 : T_809;
  assign T_812 = io_out_ready & io_out_valid;
  assign T_813 = T_812 & T_810;
  assign T_817 = T_794 + 3'h1;
  assign T_818 = T_817[2:0];
  assign GEN_175 = T_813 ? io_chosen : T_796;
  assign GEN_176 = T_813 ? T_818 : T_794;
  assign GEN_177 = T_798 ? T_796 : choice;
  assign GEN_178 = T_812 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_826 = validMask_1 | validMask_2;
  assign T_827 = T_826 | validMask_3;
  assign T_828 = T_827 | io_in_0_valid;
  assign T_829 = T_828 | io_in_1_valid;
  assign T_830 = T_829 | io_in_2_valid;
  assign T_834 = validMask_1 == 1'h0;
  assign T_836 = T_826 == 1'h0;
  assign T_838 = T_827 == 1'h0;
  assign T_840 = T_828 == 1'h0;
  assign T_842 = T_829 == 1'h0;
  assign T_844 = T_830 == 1'h0;
  assign T_848 = grantMask_1 | T_840;
  assign T_849 = T_834 & grantMask_2;
  assign T_850 = T_849 | T_842;
  assign T_851 = T_836 & grantMask_3;
  assign T_852 = T_851 | T_844;
  assign T_854 = T_796 == 2'h0;
  assign T_855 = T_798 ? T_854 : T_838;
  assign T_856 = T_855 & io_out_ready;
  assign T_858 = T_796 == 2'h1;
  assign T_859 = T_798 ? T_858 : T_848;
  assign T_860 = T_859 & io_out_ready;
  assign T_862 = T_796 == 2'h2;
  assign T_863 = T_798 ? T_862 : T_850;
  assign T_864 = T_863 & io_out_ready;
  assign T_866 = T_796 == 2'h3;
  assign T_867 = T_798 ? T_866 : T_852;
  assign T_868 = T_867 & io_out_ready;
  assign GEN_179 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_180 = io_in_1_valid ? 2'h1 : GEN_179;
  assign GEN_181 = io_in_0_valid ? 2'h0 : GEN_180;
  assign GEN_182 = validMask_3 ? 2'h3 : GEN_181;
  assign GEN_183 = validMask_2 ? 2'h2 : GEN_182;
  assign GEN_184 = validMask_1 ? 2'h1 : GEN_183;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_794 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_796 = GEN_2[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  lastGrant = GEN_3[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_794 <= 3'h0;
    end else begin
      if(T_813) begin
        T_794 <= T_818;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_813) begin
        T_796 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_812) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIORouter_1(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [10:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [10:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [10:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [10:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire [2:0] T_1855_0;
  wire [2:0] T_1855_1;
  wire  T_1857;
  wire  T_1858;
  wire  T_1859;
  wire  T_1860;
  wire [2:0] T_1861;
  wire [2:0] T_1863;
  wire [28:0] T_1864;
  wire [31:0] T_1865;
  wire  T_1869;
  wire  T_1872;
  wire  T_1874;
  wire  T_1875;
  wire  T_1877;
  wire  T_1879;
  wire  T_1880;
  wire  T_1882;
  wire  T_1884;
  wire  T_1885;
  wire [1:0] T_1886;
  wire [1:0] T_1887;
  wire [3:0] acq_route;
  wire  T_1889;
  wire  T_1890;
  wire  GEN_0;
  wire  T_1892;
  wire  T_1893;
  wire  GEN_1;
  wire  T_1895;
  wire  T_1896;
  wire  GEN_2;
  wire  T_1898;
  wire  T_1899;
  wire  GEN_3;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_2_ready;
  wire  gnt_arb_io_in_2_valid;
  wire [2:0] gnt_arb_io_in_2_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_2_bits_client_xact_id;
  wire  gnt_arb_io_in_2_bits_manager_xact_id;
  wire  gnt_arb_io_in_2_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_2_bits_g_type;
  wire [63:0] gnt_arb_io_in_2_bits_data;
  wire  gnt_arb_io_in_3_ready;
  wire  gnt_arb_io_in_3_valid;
  wire [2:0] gnt_arb_io_in_3_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_3_bits_client_xact_id;
  wire  gnt_arb_io_in_3_bits_manager_xact_id;
  wire  gnt_arb_io_in_3_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_3_bits_g_type;
  wire [63:0] gnt_arb_io_in_3_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire [1:0] gnt_arb_io_chosen;
  wire  T_1924;
  wire  T_1926;
  wire  T_1927;
  wire  T_1928;
  wire  T_1930;
  LockingRRArbiter_11 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_2_ready(gnt_arb_io_in_2_ready),
    .io_in_2_valid(gnt_arb_io_in_2_valid),
    .io_in_2_bits_addr_beat(gnt_arb_io_in_2_bits_addr_beat),
    .io_in_2_bits_client_xact_id(gnt_arb_io_in_2_bits_client_xact_id),
    .io_in_2_bits_manager_xact_id(gnt_arb_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_is_builtin_type(gnt_arb_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_g_type(gnt_arb_io_in_2_bits_g_type),
    .io_in_2_bits_data(gnt_arb_io_in_2_bits_data),
    .io_in_3_ready(gnt_arb_io_in_3_ready),
    .io_in_3_valid(gnt_arb_io_in_3_valid),
    .io_in_3_bits_addr_beat(gnt_arb_io_in_3_bits_addr_beat),
    .io_in_3_bits_client_xact_id(gnt_arb_io_in_3_bits_client_xact_id),
    .io_in_3_bits_manager_xact_id(gnt_arb_io_in_3_bits_manager_xact_id),
    .io_in_3_bits_is_builtin_type(gnt_arb_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_g_type(gnt_arb_io_in_3_bits_g_type),
    .io_in_3_bits_data(gnt_arb_io_in_3_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_3;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_1890;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign io_out_1_acquire_valid = T_1893;
  assign io_out_1_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_1_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_1_grant_ready = gnt_arb_io_in_1_ready;
  assign io_out_2_acquire_valid = T_1896;
  assign io_out_2_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_2_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_2_grant_ready = gnt_arb_io_in_2_ready;
  assign io_out_3_acquire_valid = T_1899;
  assign io_out_3_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_3_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_3_grant_ready = gnt_arb_io_in_3_ready;
  assign T_1855_0 = 3'h0;
  assign T_1855_1 = 3'h4;
  assign T_1857 = io_in_acquire_bits_a_type == T_1855_0;
  assign T_1858 = io_in_acquire_bits_a_type == T_1855_1;
  assign T_1859 = T_1857 | T_1858;
  assign T_1860 = io_in_acquire_bits_is_builtin_type & T_1859;
  assign T_1861 = io_in_acquire_bits_union[10:8];
  assign T_1863 = T_1860 ? T_1861 : 3'h0;
  assign T_1864 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_1865 = {T_1864,T_1863};
  assign T_1869 = T_1865 < 32'h1000;
  assign T_1872 = 32'h1000 <= T_1865;
  assign T_1874 = T_1865 < 32'h2000;
  assign T_1875 = T_1872 & T_1874;
  assign T_1877 = 32'h40000000 <= T_1865;
  assign T_1879 = T_1865 < 32'h44000000;
  assign T_1880 = T_1877 & T_1879;
  assign T_1882 = 32'h44000000 <= T_1865;
  assign T_1884 = T_1865 < 32'h48000000;
  assign T_1885 = T_1882 & T_1884;
  assign T_1886 = {T_1875,T_1869};
  assign T_1887 = {T_1885,T_1880};
  assign acq_route = {T_1887,T_1886};
  assign T_1889 = acq_route[0];
  assign T_1890 = io_in_acquire_valid & T_1889;
  assign GEN_0 = T_1889 ? io_out_0_acquire_ready : 1'h0;
  assign T_1892 = acq_route[1];
  assign T_1893 = io_in_acquire_valid & T_1892;
  assign GEN_1 = T_1892 ? io_out_1_acquire_ready : GEN_0;
  assign T_1895 = acq_route[2];
  assign T_1896 = io_in_acquire_valid & T_1895;
  assign GEN_2 = T_1895 ? io_out_2_acquire_ready : GEN_1;
  assign T_1898 = acq_route[3];
  assign T_1899 = io_in_acquire_valid & T_1898;
  assign GEN_3 = T_1898 ? io_out_3_acquire_ready : GEN_2;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_in_1_valid = io_out_1_grant_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = io_out_1_grant_bits_g_type;
  assign gnt_arb_io_in_1_bits_data = io_out_1_grant_bits_data;
  assign gnt_arb_io_in_2_valid = io_out_2_grant_valid;
  assign gnt_arb_io_in_2_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign gnt_arb_io_in_2_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign gnt_arb_io_in_2_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_2_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_2_bits_g_type = io_out_2_grant_bits_g_type;
  assign gnt_arb_io_in_2_bits_data = io_out_2_grant_bits_data;
  assign gnt_arb_io_in_3_valid = io_out_3_grant_valid;
  assign gnt_arb_io_in_3_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign gnt_arb_io_in_3_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign gnt_arb_io_in_3_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_3_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_3_bits_g_type = io_out_3_grant_bits_g_type;
  assign gnt_arb_io_in_3_bits_data = io_out_3_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_1924 = io_in_acquire_valid == 1'h0;
  assign T_1926 = acq_route != 4'h0;
  assign T_1927 = T_1924 | T_1926;
  assign T_1928 = T_1927 | reset;
  assign T_1930 = T_1928 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1930) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at Interconnect.scala:219 assert(!io.in.acquire.valid || acq_route.orR, \"No valid route\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1930) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [10:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [10:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [10:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_1_1_clk;
  wire  ClientUncachedTileLinkIORouter_1_1_reset;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data;
  ClientUncachedTileLinkIORouter_1 ClientUncachedTileLinkIORouter_1_1 (
    .clk(ClientUncachedTileLinkIORouter_1_1_clk),
    .reset(ClientUncachedTileLinkIORouter_1_1_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready),
    .io_out_2_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready),
    .io_out_3_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_1_clk = clk;
  assign ClientUncachedTileLinkIORouter_1_1_reset = reset;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid = io_out_2_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid = io_out_3_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [10:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [10:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [10:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [10:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [10:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  xbar_io_out_1_acquire_ready;
  wire  xbar_io_out_1_acquire_valid;
  wire [25:0] xbar_io_out_1_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_1_acquire_bits_addr_beat;
  wire  xbar_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_1_acquire_bits_a_type;
  wire [10:0] xbar_io_out_1_acquire_bits_union;
  wire [63:0] xbar_io_out_1_acquire_bits_data;
  wire  xbar_io_out_1_grant_ready;
  wire  xbar_io_out_1_grant_valid;
  wire [2:0] xbar_io_out_1_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_1_grant_bits_client_xact_id;
  wire  xbar_io_out_1_grant_bits_manager_xact_id;
  wire  xbar_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_1_grant_bits_g_type;
  wire [63:0] xbar_io_out_1_grant_bits_data;
  wire  xbar_io_out_2_acquire_ready;
  wire  xbar_io_out_2_acquire_valid;
  wire [25:0] xbar_io_out_2_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_2_acquire_bits_addr_beat;
  wire  xbar_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_2_acquire_bits_a_type;
  wire [10:0] xbar_io_out_2_acquire_bits_union;
  wire [63:0] xbar_io_out_2_acquire_bits_data;
  wire  xbar_io_out_2_grant_ready;
  wire  xbar_io_out_2_grant_valid;
  wire [2:0] xbar_io_out_2_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_2_grant_bits_client_xact_id;
  wire  xbar_io_out_2_grant_bits_manager_xact_id;
  wire  xbar_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_2_grant_bits_g_type;
  wire [63:0] xbar_io_out_2_grant_bits_data;
  wire  xbar_io_out_3_acquire_ready;
  wire  xbar_io_out_3_acquire_valid;
  wire [25:0] xbar_io_out_3_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_3_acquire_bits_addr_beat;
  wire  xbar_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_3_acquire_bits_a_type;
  wire [10:0] xbar_io_out_3_acquire_bits_union;
  wire [63:0] xbar_io_out_3_acquire_bits_data;
  wire  xbar_io_out_3_grant_ready;
  wire  xbar_io_out_3_grant_valid;
  wire [2:0] xbar_io_out_3_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_3_grant_bits_client_xact_id;
  wire  xbar_io_out_3_grant_bits_manager_xact_id;
  wire  xbar_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_3_grant_bits_g_type;
  wire [63:0] xbar_io_out_3_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar_1 xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(xbar_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(xbar_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(xbar_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(xbar_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(xbar_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(xbar_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(xbar_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(xbar_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(xbar_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(xbar_io_out_1_grant_ready),
    .io_out_1_grant_valid(xbar_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(xbar_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(xbar_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(xbar_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(xbar_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(xbar_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(xbar_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(xbar_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(xbar_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(xbar_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(xbar_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(xbar_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(xbar_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(xbar_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(xbar_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(xbar_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(xbar_io_out_2_grant_ready),
    .io_out_2_grant_valid(xbar_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(xbar_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(xbar_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(xbar_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(xbar_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(xbar_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(xbar_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(xbar_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(xbar_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(xbar_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(xbar_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(xbar_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(xbar_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(xbar_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(xbar_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(xbar_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(xbar_io_out_3_grant_ready),
    .io_out_3_grant_valid(xbar_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(xbar_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(xbar_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(xbar_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(xbar_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(xbar_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(xbar_io_out_3_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = xbar_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = xbar_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = xbar_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = xbar_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = xbar_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = xbar_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = xbar_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = xbar_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = xbar_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = xbar_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = xbar_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = xbar_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = xbar_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = xbar_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = xbar_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = xbar_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = xbar_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = xbar_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = xbar_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = xbar_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = xbar_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = xbar_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = xbar_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = xbar_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = xbar_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = xbar_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = xbar_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = xbar_io_out_3_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = io_out_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign xbar_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign xbar_io_out_1_grant_valid = io_out_1_grant_valid;
  assign xbar_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign xbar_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign xbar_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign xbar_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign xbar_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign xbar_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign xbar_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign xbar_io_out_2_grant_valid = io_out_2_grant_valid;
  assign xbar_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign xbar_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign xbar_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign xbar_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign xbar_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign xbar_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign xbar_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign xbar_io_out_3_grant_valid = io_out_3_grant_valid;
  assign xbar_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign xbar_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign xbar_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign xbar_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign xbar_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign xbar_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [10:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [10:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [10:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [10:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [10:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_clk;
  wire  TileLinkRecursiveInterconnect_1_1_reset;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data)
  );
  TileLinkRecursiveInterconnect_1 TileLinkRecursiveInterconnect_1_1 (
    .clk(TileLinkRecursiveInterconnect_1_1_clk),
    .reset(TileLinkRecursiveInterconnect_1_1_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_clk = clk;
  assign TileLinkRecursiveInterconnect_1_1_reset = reset;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready = xbar_io_out_0_grant_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid = io_out_2_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid = io_out_3_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
endmodule
module Queue_12(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [25:0] io_enq_bits_addr_block,
  input  [1:0] io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input  [10:0] io_enq_bits_union,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [25:0] io_deq_bits_addr_block,
  output [1:0] io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [10:0] io_deq_bits_union,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [25:0] ram_addr_block [0:0];
  reg [31:0] GEN_0;
  wire [25:0] ram_addr_block_T_254_data;
  wire  ram_addr_block_T_254_addr;
  wire  ram_addr_block_T_254_en;
  wire [25:0] ram_addr_block_T_224_data;
  wire  ram_addr_block_T_224_addr;
  wire  ram_addr_block_T_224_mask;
  wire  ram_addr_block_T_224_en;
  reg [1:0] ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_client_xact_id_T_254_data;
  wire  ram_client_xact_id_T_254_addr;
  wire  ram_client_xact_id_T_254_en;
  wire [1:0] ram_client_xact_id_T_224_data;
  wire  ram_client_xact_id_T_224_addr;
  wire  ram_client_xact_id_T_224_mask;
  wire  ram_client_xact_id_T_224_en;
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_addr_beat_T_254_data;
  wire  ram_addr_beat_T_254_addr;
  wire  ram_addr_beat_T_254_en;
  wire [2:0] ram_addr_beat_T_224_data;
  wire  ram_addr_beat_T_224_addr;
  wire  ram_addr_beat_T_224_mask;
  wire  ram_addr_beat_T_224_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_254_data;
  wire  ram_is_builtin_type_T_254_addr;
  wire  ram_is_builtin_type_T_254_en;
  wire  ram_is_builtin_type_T_224_data;
  wire  ram_is_builtin_type_T_224_addr;
  wire  ram_is_builtin_type_T_224_mask;
  wire  ram_is_builtin_type_T_224_en;
  reg [2:0] ram_a_type [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_254_data;
  wire  ram_a_type_T_254_addr;
  wire  ram_a_type_T_254_en;
  wire [2:0] ram_a_type_T_224_data;
  wire  ram_a_type_T_224_addr;
  wire  ram_a_type_T_224_mask;
  wire  ram_a_type_T_224_en;
  reg [10:0] ram_union [0:0];
  reg [31:0] GEN_5;
  wire [10:0] ram_union_T_254_data;
  wire  ram_union_T_254_addr;
  wire  ram_union_T_254_en;
  wire [10:0] ram_union_T_224_data;
  wire  ram_union_T_224_addr;
  wire  ram_union_T_224_mask;
  wire  ram_union_T_224_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_6;
  wire [63:0] ram_data_T_254_data;
  wire  ram_data_T_254_addr;
  wire  ram_data_T_254_en;
  wire [63:0] ram_data_T_224_data;
  wire  ram_data_T_224_addr;
  wire  ram_data_T_224_mask;
  wire  ram_data_T_224_en;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  T_221;
  wire  T_222;
  wire  do_enq;
  wire  T_223;
  wire  do_deq;
  wire  T_249;
  wire  GEN_17;
  wire  T_251;
  wire [1:0] T_277;
  wire  ptr_diff;
  wire [1:0] T_279;
  assign io_enq_ready = T_221;
  assign io_deq_valid = T_251;
  assign io_deq_bits_addr_block = ram_addr_block_T_254_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_254_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_254_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_254_data;
  assign io_deq_bits_a_type = ram_a_type_T_254_data;
  assign io_deq_bits_union = ram_union_T_254_data;
  assign io_deq_bits_data = ram_data_T_254_data;
  assign io_count = T_279[0];
  assign ram_addr_block_T_254_addr = 1'h0;
  assign ram_addr_block_T_254_en = 1'h1;
  assign ram_addr_block_T_254_data = ram_addr_block[ram_addr_block_T_254_addr];
  assign ram_addr_block_T_224_data = io_enq_bits_addr_block;
  assign ram_addr_block_T_224_addr = 1'h0;
  assign ram_addr_block_T_224_mask = do_enq;
  assign ram_addr_block_T_224_en = do_enq;
  assign ram_client_xact_id_T_254_addr = 1'h0;
  assign ram_client_xact_id_T_254_en = 1'h1;
  assign ram_client_xact_id_T_254_data = ram_client_xact_id[ram_client_xact_id_T_254_addr];
  assign ram_client_xact_id_T_224_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_224_addr = 1'h0;
  assign ram_client_xact_id_T_224_mask = do_enq;
  assign ram_client_xact_id_T_224_en = do_enq;
  assign ram_addr_beat_T_254_addr = 1'h0;
  assign ram_addr_beat_T_254_en = 1'h1;
  assign ram_addr_beat_T_254_data = ram_addr_beat[ram_addr_beat_T_254_addr];
  assign ram_addr_beat_T_224_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_224_addr = 1'h0;
  assign ram_addr_beat_T_224_mask = do_enq;
  assign ram_addr_beat_T_224_en = do_enq;
  assign ram_is_builtin_type_T_254_addr = 1'h0;
  assign ram_is_builtin_type_T_254_en = 1'h1;
  assign ram_is_builtin_type_T_254_data = ram_is_builtin_type[ram_is_builtin_type_T_254_addr];
  assign ram_is_builtin_type_T_224_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_224_addr = 1'h0;
  assign ram_is_builtin_type_T_224_mask = do_enq;
  assign ram_is_builtin_type_T_224_en = do_enq;
  assign ram_a_type_T_254_addr = 1'h0;
  assign ram_a_type_T_254_en = 1'h1;
  assign ram_a_type_T_254_data = ram_a_type[ram_a_type_T_254_addr];
  assign ram_a_type_T_224_data = io_enq_bits_a_type;
  assign ram_a_type_T_224_addr = 1'h0;
  assign ram_a_type_T_224_mask = do_enq;
  assign ram_a_type_T_224_en = do_enq;
  assign ram_union_T_254_addr = 1'h0;
  assign ram_union_T_254_en = 1'h1;
  assign ram_union_T_254_data = ram_union[ram_union_T_254_addr];
  assign ram_union_T_224_data = io_enq_bits_union;
  assign ram_union_T_224_addr = 1'h0;
  assign ram_union_T_224_mask = do_enq;
  assign ram_union_T_224_en = do_enq;
  assign ram_data_T_254_addr = 1'h0;
  assign ram_data_T_254_en = 1'h1;
  assign ram_data_T_254_data = ram_data[ram_data_T_254_addr];
  assign ram_data_T_224_data = io_enq_bits_data;
  assign ram_data_T_224_addr = 1'h0;
  assign ram_data_T_224_mask = do_enq;
  assign ram_data_T_224_en = do_enq;
  assign T_221 = maybe_full == 1'h0;
  assign T_222 = io_enq_ready & io_enq_valid;
  assign do_enq = T_222;
  assign T_223 = io_deq_ready & io_deq_valid;
  assign do_deq = T_223;
  assign T_249 = do_enq != do_deq;
  assign GEN_17 = T_249 ? do_enq : maybe_full;
  assign T_251 = T_221 == 1'h0;
  assign T_277 = 1'h0 - 1'h0;
  assign ptr_diff = T_277[0:0];
  assign T_279 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_block[initvar] = GEN_0[25:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_union[initvar] = GEN_5[10:0];
  `endif
  GEN_6 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_6[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_block_T_224_en & ram_addr_block_T_224_mask) begin
      ram_addr_block[ram_addr_block_T_224_addr] <= ram_addr_block_T_224_data;
    end
    if(ram_client_xact_id_T_224_en & ram_client_xact_id_T_224_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_224_addr] <= ram_client_xact_id_T_224_data;
    end
    if(ram_addr_beat_T_224_en & ram_addr_beat_T_224_mask) begin
      ram_addr_beat[ram_addr_beat_T_224_addr] <= ram_addr_beat_T_224_data;
    end
    if(ram_is_builtin_type_T_224_en & ram_is_builtin_type_T_224_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_224_addr] <= ram_is_builtin_type_T_224_data;
    end
    if(ram_a_type_T_224_en & ram_a_type_T_224_mask) begin
      ram_a_type[ram_a_type_T_224_addr] <= ram_a_type_T_224_data;
    end
    if(ram_union_T_224_en & ram_union_T_224_mask) begin
      ram_union[ram_union_T_224_addr] <= ram_union_T_224_data;
    end
    if(ram_data_T_224_en & ram_data_T_224_mask) begin
      ram_data[ram_data_T_224_addr] <= ram_data_T_224_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_249) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module PLIC(
  input   clk,
  input   reset,
  input   io_devices_0_valid,
  output  io_devices_0_ready,
  output  io_devices_0_complete,
  input   io_devices_1_valid,
  output  io_devices_1_ready,
  output  io_devices_1_complete,
  output  io_harts_0,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [10:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data
);
  wire  T_477_0;
  wire  T_477_1;
  wire  T_477_2;
  wire  priority_0;
  wire  priority_1;
  wire  priority_2;
  wire  T_488_0;
  wire  threshold_0;
  wire  T_501_0;
  wire  T_501_1;
  wire  T_501_2;
  reg  pending_0;
  reg [31:0] GEN_8;
  reg  pending_1;
  reg [31:0] GEN_14;
  reg  pending_2;
  reg [31:0] GEN_17;
  reg  enables_0_0;
  reg [31:0] GEN_18;
  reg  enables_0_1;
  reg [31:0] GEN_19;
  reg  enables_0_2;
  reg [31:0] GEN_26;
  wire  T_538;
  wire  GEN_12;
  wire  T_542;
  wire  GEN_13;
  wire [1:0] maxDevs_0;
  wire  T_552;
  wire [1:0] T_553;
  wire  T_554;
  wire [1:0] T_555;
  wire  T_560;
  wire [1:0] T_561;
  wire [1:0] T_563;
  wire  T_564;
  wire  T_565;
  wire  T_567;
  wire [1:0] T_568;
  wire [2:0] T_570;
  wire [1:0] T_571;
  wire [1:0] T_572;
  reg [1:0] T_573;
  reg [31:0] GEN_29;
  reg [1:0] T_574;
  reg [31:0] GEN_30;
  wire [1:0] T_576;
  wire  T_577;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [10:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [10:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_601;
  wire  T_603;
  wire  T_604;
  wire  read;
  wire  T_607;
  wire  T_608;
  wire  write;
  wire  T_611;
  wire  T_612;
  wire  T_613;
  wire  T_614;
  wire  T_616;
  wire [2:0] T_624_0;
  wire [2:0] T_624_1;
  wire  T_626;
  wire  T_627;
  wire  T_628;
  wire  T_629;
  wire [2:0] T_630;
  wire [2:0] T_632;
  wire [28:0] T_633;
  wire [31:0] T_634;
  wire [25:0] addr;
  wire  hart;
  wire [63:0] rdata;
  wire  T_640;
  wire  T_641;
  wire  T_660;
  wire  T_661;
  wire  T_665;
  wire [7:0] T_666;
  wire [7:0] T_668;
  wire [7:0] T_669;
  wire  T_670;
  wire  T_671;
  wire  T_672;
  wire  T_673;
  wire  T_674;
  wire  T_675;
  wire  T_676;
  wire  T_677;
  wire [7:0] T_681;
  wire [7:0] T_685;
  wire [7:0] T_689;
  wire [7:0] T_693;
  wire [7:0] T_697;
  wire [7:0] T_701;
  wire [7:0] T_705;
  wire [7:0] T_709;
  wire [15:0] T_710;
  wire [15:0] T_711;
  wire [31:0] T_712;
  wire [15:0] T_713;
  wire [15:0] T_714;
  wire [31:0] T_715;
  wire [63:0] T_716;
  wire [63:0] T_717;
  wire [63:0] T_796;
  wire [63:0] T_797;
  wire [63:0] masked_wdata;
  wire  T_799;
  wire [1:0] GEN_0;
  wire [32:0] T_802;
  wire  GEN_1;
  wire [33:0] T_803;
  wire [7:0] T_805;
  wire [33:0] T_806;
  wire  T_807;
  wire  T_808;
  wire [1:0] GEN_2;
  wire  GEN_3;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_20;
  wire  GEN_21;
  wire [31:0] T_842;
  wire [1:0] T_843;
  wire  GEN_4;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_22;
  wire  GEN_95;
  wire  GEN_23;
  wire [2:0] T_845;
  wire [1:0] T_846;
  wire  GEN_5;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_35;
  wire  GEN_36;
  wire [63:0] GEN_39;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_47;
  wire  GEN_48;
  wire  T_854;
  wire  T_856;
  wire  T_857;
  wire  GEN_6_0;
  wire  GEN_6_1;
  wire  GEN_6_2;
  wire  GEN_7_0;
  wire  GEN_7_1;
  wire  GEN_7_2;
  wire [1:0] T_862;
  wire  GEN_8_0;
  wire  GEN_8_1;
  wire  GEN_8_2;
  wire [2:0] T_863;
  wire  T_867;
  wire  GEN_9;
  wire  T_871;
  wire  GEN_10;
  wire  GEN_54;
  wire  T_875;
  wire  GEN_11;
  wire  GEN_57;
  wire [63:0] GEN_67;
  wire [63:0] GEN_84;
  wire  GEN_88;
  wire  GEN_90;
  wire  T_877;
  wire  T_881;
  wire  T_882;
  wire  T_883;
  wire [1:0] T_885;
  wire [2:0] T_886;
  wire [2:0] T_889;
  wire [63:0] GEN_91;
  wire  T_896;
  wire  T_897;
  wire  T_898;
  wire  T_900;
  wire [31:0] T_902;
  wire [31:0] T_904;
  wire [63:0] T_905;
  wire [63:0] GEN_92;
  wire [31:0] T_909;
  wire [63:0] GEN_93;
  wire [63:0] GEN_94;
  wire  T_929;
  wire [2:0] T_930;
  wire  T_931;
  wire [2:0] T_932;
  wire  T_933;
  wire [2:0] T_934;
  wire  T_935;
  wire [2:0] T_936;
  wire  T_937;
  wire [2:0] T_938;
  wire  T_939;
  wire [2:0] T_940;
  wire  T_941;
  wire [2:0] T_942;
  wire [2:0] T_967_addr_beat;
  wire [1:0] T_967_client_xact_id;
  wire  T_967_manager_xact_id;
  wire  T_967_is_builtin_type;
  wire [3:0] T_967_g_type;
  wire [63:0] T_967_data;
  Queue_12 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_devices_0_ready = T_538;
  assign io_devices_0_complete = GEN_47;
  assign io_devices_1_ready = T_542;
  assign io_devices_1_complete = GEN_48;
  assign io_harts_0 = T_577;
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_967_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_967_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_967_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_967_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_967_g_type;
  assign io_tl_grant_bits_data = T_967_data;
  assign T_477_0 = 1'h1;
  assign T_477_1 = 1'h1;
  assign T_477_2 = 1'h1;
  assign priority_0 = 1'h0;
  assign priority_1 = T_477_1;
  assign priority_2 = T_477_2;
  assign T_488_0 = 1'h0;
  assign threshold_0 = T_488_0;
  assign T_501_0 = 1'h0;
  assign T_501_1 = 1'h0;
  assign T_501_2 = 1'h0;
  assign T_538 = pending_1 == 1'h0;
  assign GEN_12 = io_devices_0_valid ? 1'h1 : pending_1;
  assign T_542 = pending_2 == 1'h0;
  assign GEN_13 = io_devices_1_valid ? 1'h1 : pending_2;
  assign maxDevs_0 = T_573;
  assign T_552 = pending_1 & enables_0_1;
  assign T_553 = {T_552,priority_1};
  assign T_554 = pending_2 & enables_0_2;
  assign T_555 = {T_554,priority_2};
  assign T_560 = 2'h2 >= T_553;
  assign T_561 = T_560 ? 2'h2 : T_553;
  assign T_563 = 1'h1 + 1'h0;
  assign T_564 = T_563[0:0];
  assign T_565 = T_560 ? 1'h0 : T_564;
  assign T_567 = T_561 >= T_555;
  assign T_568 = T_567 ? T_561 : T_555;
  assign T_570 = 2'h2 + 2'h0;
  assign T_571 = T_570[1:0];
  assign T_572 = T_567 ? {{1'd0}, T_565} : T_571;
  assign T_576 = {1'h1,threshold_0};
  assign T_577 = T_574 > T_576;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_601 = acq_io_deq_ready & acq_io_deq_valid;
  assign T_603 = acq_io_deq_bits_a_type == 3'h0;
  assign T_604 = acq_io_deq_bits_is_builtin_type & T_603;
  assign read = T_601 & T_604;
  assign T_607 = acq_io_deq_bits_a_type == 3'h2;
  assign T_608 = acq_io_deq_bits_is_builtin_type & T_607;
  assign write = T_601 & T_608;
  assign T_611 = T_601 == 1'h0;
  assign T_612 = T_611 | read;
  assign T_613 = T_612 | write;
  assign T_614 = T_613 | reset;
  assign T_616 = T_614 == 1'h0;
  assign T_624_0 = 3'h0;
  assign T_624_1 = 3'h4;
  assign T_626 = acq_io_deq_bits_a_type == T_624_0;
  assign T_627 = acq_io_deq_bits_a_type == T_624_1;
  assign T_628 = T_626 | T_627;
  assign T_629 = acq_io_deq_bits_is_builtin_type & T_628;
  assign T_630 = acq_io_deq_bits_union[10:8];
  assign T_632 = T_629 ? T_630 : 3'h0;
  assign T_633 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_634 = {T_633,T_632};
  assign addr = T_634[25:0];
  assign hart = 1'h0;
  assign rdata = GEN_94;
  assign T_640 = acq_io_deq_bits_a_type == 3'h4;
  assign T_641 = acq_io_deq_bits_is_builtin_type & T_640;
  assign T_660 = acq_io_deq_bits_a_type == 3'h3;
  assign T_661 = acq_io_deq_bits_is_builtin_type & T_660;
  assign T_665 = T_661 | T_608;
  assign T_666 = acq_io_deq_bits_union[8:1];
  assign T_668 = T_665 ? T_666 : 8'h0;
  assign T_669 = T_641 ? 8'hff : T_668;
  assign T_670 = T_669[0];
  assign T_671 = T_669[1];
  assign T_672 = T_669[2];
  assign T_673 = T_669[3];
  assign T_674 = T_669[4];
  assign T_675 = T_669[5];
  assign T_676 = T_669[6];
  assign T_677 = T_669[7];
  assign T_681 = T_670 ? 8'hff : 8'h0;
  assign T_685 = T_671 ? 8'hff : 8'h0;
  assign T_689 = T_672 ? 8'hff : 8'h0;
  assign T_693 = T_673 ? 8'hff : 8'h0;
  assign T_697 = T_674 ? 8'hff : 8'h0;
  assign T_701 = T_675 ? 8'hff : 8'h0;
  assign T_705 = T_676 ? 8'hff : 8'h0;
  assign T_709 = T_677 ? 8'hff : 8'h0;
  assign T_710 = {T_685,T_681};
  assign T_711 = {T_693,T_689};
  assign T_712 = {T_711,T_710};
  assign T_713 = {T_701,T_697};
  assign T_714 = {T_709,T_705};
  assign T_715 = {T_714,T_713};
  assign T_716 = {T_715,T_712};
  assign T_717 = acq_io_deq_bits_data & T_716;
  assign T_796 = ~ T_716;
  assign T_797 = rdata & T_796;
  assign masked_wdata = T_717 | T_797;
  assign T_799 = addr >= 26'h200000;
  assign GEN_0 = maxDevs_0;
  assign T_802 = {GEN_0,31'h0};
  assign GEN_1 = threshold_0;
  assign T_803 = {T_802,GEN_1};
  assign T_805 = 7'h0 * 7'h40;
  assign T_806 = T_803 >> T_805;
  assign T_807 = addr[2];
  assign T_808 = read & T_807;
  assign GEN_2 = maxDevs_0;
  assign GEN_3 = 1'h0;
  assign GEN_15 = 2'h1 == GEN_2 ? GEN_3 : GEN_12;
  assign GEN_16 = 2'h2 == GEN_2 ? GEN_3 : GEN_13;
  assign GEN_20 = T_808 ? GEN_15 : GEN_12;
  assign GEN_21 = T_808 ? GEN_16 : GEN_13;
  assign T_842 = acq_io_deq_bits_data[63:32];
  assign T_843 = T_842[1:0];
  assign GEN_4 = GEN_23;
  assign GEN_6 = 1'h0 == hart;
  assign GEN_7 = 2'h1 == T_843;
  assign GEN_22 = GEN_6 & GEN_7 ? enables_0_1 : enables_0_0;
  assign GEN_95 = 2'h2 == T_843;
  assign GEN_23 = GEN_6 & GEN_95 ? enables_0_2 : GEN_22;
  assign T_845 = T_843 - 2'h1;
  assign T_846 = T_845[1:0];
  assign GEN_5 = 1'h1;
  assign GEN_24 = 2'h0 == T_846 ? GEN_5 : 1'h0;
  assign GEN_25 = 2'h1 == T_846 ? GEN_5 : 1'h0;
  assign GEN_27 = GEN_4 ? GEN_24 : 1'h0;
  assign GEN_28 = GEN_4 ? GEN_25 : 1'h0;
  assign GEN_31 = T_674 ? GEN_27 : 1'h0;
  assign GEN_32 = T_674 ? GEN_28 : 1'h0;
  assign GEN_35 = write ? GEN_31 : 1'h0;
  assign GEN_36 = write ? GEN_32 : 1'h0;
  assign GEN_39 = T_799 ? {{30'd0}, T_806} : 64'h0;
  assign GEN_43 = T_799 ? GEN_20 : GEN_12;
  assign GEN_44 = T_799 ? GEN_21 : GEN_13;
  assign GEN_47 = T_799 ? GEN_35 : 1'h0;
  assign GEN_48 = T_799 ? GEN_36 : 1'h0;
  assign T_854 = addr >= 26'h2000;
  assign T_856 = T_799 == 1'h0;
  assign T_857 = T_856 & T_854;
  assign GEN_6_0 = enables_0_0;
  assign GEN_6_1 = enables_0_1;
  assign GEN_6_2 = enables_0_2;
  assign GEN_7_0 = enables_0_0;
  assign GEN_7_1 = enables_0_1;
  assign GEN_7_2 = enables_0_2;
  assign T_862 = {GEN_6_2,GEN_7_1};
  assign GEN_8_0 = enables_0_0;
  assign GEN_8_1 = enables_0_1;
  assign GEN_8_2 = enables_0_2;
  assign T_863 = {T_862,GEN_8_0};
  assign T_867 = masked_wdata[0];
  assign GEN_9 = T_867;
  assign T_871 = masked_wdata[1];
  assign GEN_10 = T_871;
  assign GEN_54 = write ? GEN_10 : enables_0_1;
  assign T_875 = masked_wdata[2];
  assign GEN_11 = T_875;
  assign GEN_57 = write ? GEN_11 : enables_0_2;
  assign GEN_67 = {{61'd0}, T_863};
  assign GEN_84 = T_857 ? GEN_67 : GEN_39;
  assign GEN_88 = T_857 ? GEN_54 : enables_0_1;
  assign GEN_90 = T_857 ? GEN_57 : enables_0_2;
  assign T_877 = addr >= 26'h1000;
  assign T_881 = T_854 == 1'h0;
  assign T_882 = T_856 & T_881;
  assign T_883 = T_882 & T_877;
  assign T_885 = {pending_2,pending_1};
  assign T_886 = {T_885,pending_0};
  assign T_889 = T_886 >> T_805;
  assign GEN_91 = T_883 ? {{61'd0}, T_889} : GEN_84;
  assign T_896 = T_877 == 1'h0;
  assign T_897 = T_882 & T_896;
  assign T_898 = addr[3];
  assign T_900 = T_898 == 1'h0;
  assign T_902 = {31'h0,priority_0};
  assign T_904 = {31'h0,priority_1};
  assign T_905 = {T_904,T_902};
  assign GEN_92 = T_900 ? T_905 : GEN_91;
  assign T_909 = {31'h0,priority_2};
  assign GEN_93 = T_898 ? {{32'd0}, T_909} : GEN_92;
  assign GEN_94 = T_897 ? GEN_93 : GEN_91;
  assign T_929 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_930 = T_929 ? 3'h1 : 3'h3;
  assign T_931 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_932 = T_931 ? 3'h1 : T_930;
  assign T_933 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_934 = T_933 ? 3'h4 : T_932;
  assign T_935 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_936 = T_935 ? 3'h3 : T_934;
  assign T_937 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_938 = T_937 ? 3'h3 : T_936;
  assign T_939 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_940 = T_939 ? 3'h5 : T_938;
  assign T_941 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_942 = T_941 ? 3'h4 : T_940;
  assign T_967_addr_beat = 3'h0;
  assign T_967_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_967_manager_xact_id = 1'h0;
  assign T_967_is_builtin_type = 1'h1;
  assign T_967_g_type = {{1'd0}, T_942};
  assign T_967_data = rdata;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  pending_0 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_14 = {1{$random}};
  pending_1 = GEN_14[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {1{$random}};
  pending_2 = GEN_17[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {1{$random}};
  enables_0_0 = GEN_18[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_19 = {1{$random}};
  enables_0_1 = GEN_19[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_26 = {1{$random}};
  enables_0_2 = GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  T_573 = GEN_29[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  T_574 = GEN_30[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      pending_0 <= T_501_0;
    end else begin
      pending_0 <= 1'h0;
    end
    if(reset) begin
      pending_1 <= T_501_1;
    end else begin
      if(T_799) begin
        if(T_808) begin
          if(2'h1 == GEN_2) begin
            pending_1 <= GEN_3;
          end else begin
            if(io_devices_0_valid) begin
              pending_1 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_0_valid) begin
            pending_1 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_0_valid) begin
          pending_1 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_2 <= T_501_2;
    end else begin
      if(T_799) begin
        if(T_808) begin
          if(2'h2 == GEN_2) begin
            pending_2 <= GEN_3;
          end else begin
            if(io_devices_1_valid) begin
              pending_2 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_1_valid) begin
            pending_2 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_1_valid) begin
          pending_2 <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      enables_0_0 <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(T_857) begin
        if(write) begin
          enables_0_1 <= GEN_10;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_857) begin
        if(write) begin
          enables_0_2 <= GEN_11;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_567) begin
        T_573 <= {{1'd0}, T_565};
      end else begin
        T_573 <= T_571;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_567) begin
        if(T_560) begin
          T_574 <= 2'h2;
        end else begin
          T_574 <= T_553;
        end
      end else begin
        T_574 <= T_555;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_616) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported PLIC operation\n    at Plic.scala:108 assert(!acq.fire() || read || write, \"unsupported PLIC operation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_616) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module LevelGateway(
  input   clk,
  input   reset,
  input   io_interrupt,
  output  io_plic_valid,
  input   io_plic_ready,
  input   io_plic_complete
);
  reg  inFlight;
  reg [31:0] GEN_2;
  wire  T_6;
  wire  GEN_0;
  wire  GEN_1;
  wire  T_10;
  wire  T_11;
  assign io_plic_valid = T_11;
  assign T_6 = io_interrupt & io_plic_ready;
  assign GEN_0 = T_6 ? 1'h1 : inFlight;
  assign GEN_1 = io_plic_complete ? 1'h0 : GEN_0;
  assign T_10 = inFlight == 1'h0;
  assign T_11 = io_interrupt & T_10;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  inFlight = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      inFlight <= 1'h0;
    end else begin
      if(io_plic_complete) begin
        inFlight <= 1'h0;
      end else begin
        if(T_6) begin
          inFlight <= 1'h1;
        end
      end
    end
  end
endmodule
module DebugModule(
  input   clk,
  input   reset,
  output  io_db_req_ready,
  input   io_db_req_valid,
  input  [4:0] io_db_req_bits_addr,
  input  [33:0] io_db_req_bits_data,
  input  [1:0] io_db_req_bits_op,
  input   io_db_resp_ready,
  output  io_db_resp_valid,
  output [33:0] io_db_resp_bits_data,
  output [1:0] io_db_resp_bits_resp,
  output  io_debugInterrupts_0,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [10:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_ndreset,
  output  io_fullreset
);
  wire  CONTROLReset_interrupt;
  wire  CONTROLReset_haltnot;
  wire [9:0] CONTROLReset_reserved0;
  wire [2:0] CONTROLReset_buserror;
  wire [2:0] CONTROLReset_serial;
  wire  CONTROLReset_autoincrement;
  wire [2:0] CONTROLReset_access;
  wire [9:0] CONTROLReset_hartid;
  wire  CONTROLReset_ndreset;
  wire  CONTROLReset_fullreset;
  wire  CONTROLWrEn;
  reg  CONTROLReg_interrupt;
  reg [31:0] GEN_26;
  reg  CONTROLReg_haltnot;
  reg [31:0] GEN_27;
  reg [9:0] CONTROLReg_reserved0;
  reg [31:0] GEN_28;
  reg [2:0] CONTROLReg_buserror;
  reg [31:0] GEN_29;
  reg [2:0] CONTROLReg_serial;
  reg [31:0] GEN_30;
  reg  CONTROLReg_autoincrement;
  reg [31:0] GEN_52;
  reg [2:0] CONTROLReg_access;
  reg [31:0] GEN_85;
  reg [9:0] CONTROLReg_hartid;
  reg [31:0] GEN_86;
  reg  CONTROLReg_ndreset;
  reg [31:0] GEN_88;
  reg  CONTROLReg_fullreset;
  reg [31:0] GEN_89;
  wire  CONTROLWrData_interrupt;
  wire  CONTROLWrData_haltnot;
  wire [9:0] CONTROLWrData_reserved0;
  wire [2:0] CONTROLWrData_buserror;
  wire [2:0] CONTROLWrData_serial;
  wire  CONTROLWrData_autoincrement;
  wire [2:0] CONTROLWrData_access;
  wire [9:0] CONTROLWrData_hartid;
  wire  CONTROLWrData_ndreset;
  wire  CONTROLWrData_fullreset;
  wire  CONTROLRdData_interrupt;
  wire  CONTROLRdData_haltnot;
  wire [9:0] CONTROLRdData_reserved0;
  wire [2:0] CONTROLRdData_buserror;
  wire [2:0] CONTROLRdData_serial;
  wire  CONTROLRdData_autoincrement;
  wire [2:0] CONTROLRdData_access;
  wire [9:0] CONTROLRdData_hartid;
  wire  CONTROLRdData_ndreset;
  wire  CONTROLRdData_fullreset;
  reg  ndresetCtrReg;
  reg [31:0] GEN_90;
  wire [1:0] DMINFORdData_reserved0;
  wire [6:0] DMINFORdData_abussize;
  wire [3:0] DMINFORdData_serialcount;
  wire  DMINFORdData_access128;
  wire  DMINFORdData_access64;
  wire  DMINFORdData_access32;
  wire  DMINFORdData_access16;
  wire  DMINFORdData_accesss8;
  wire [5:0] DMINFORdData_dramsize;
  wire  DMINFORdData_haltsum;
  wire [2:0] DMINFORdData_reserved1;
  wire  DMINFORdData_authenticated;
  wire  DMINFORdData_authbusy;
  wire [1:0] DMINFORdData_authtype;
  wire [1:0] DMINFORdData_version;
  wire  HALTSUMRdData_serialfull;
  wire  HALTSUMRdData_serialvalid;
  wire [31:0] HALTSUMRdData_acks;
  wire  RAMWrData_interrupt;
  wire  RAMWrData_haltnot;
  wire [31:0] RAMWrData_data;
  wire  RAMRdData_interrupt;
  wire  RAMRdData_haltnot;
  wire [31:0] RAMRdData_data;
  wire  SETHALTNOTWrEn;
  wire [9:0] SETHALTNOTWrData;
  wire  CLEARDEBINTWrEn;
  wire [9:0] CLEARDEBINTWrData;
  wire  T_655_0;
  reg  interruptRegs_0;
  reg [31:0] GEN_109;
  wire  T_666_0;
  reg  haltnotRegs_0;
  reg [31:0] GEN_110;
  wire [31:0] haltnotStatus_0;
  wire [31:0] rdHaltnotStatus;
  wire  haltnotSummary;
  reg [63:0] ramMem [0:7];
  reg [63:0] GEN_111;
  wire [63:0] ramMem_T_850_data;
  wire [2:0] ramMem_T_850_addr;
  wire  ramMem_T_850_en;
  wire [63:0] ramMem_T_851_data;
  wire [2:0] ramMem_T_851_addr;
  wire  ramMem_T_851_mask;
  wire  ramMem_T_851_en;
  wire [2:0] ramAddr;
  wire [63:0] ramRdData;
  wire [63:0] ramWrData;
  wire [63:0] ramWrMask;
  wire  ramWrEn;
  wire [3:0] dbRamAddr;
  wire [31:0] dbRamRdData;
  wire [31:0] dbRamWrData;
  wire  dbRamWrEn;
  wire  dbRamRdEn;
  wire [2:0] sbRamAddr;
  wire [63:0] sbRamRdData;
  wire [63:0] sbRamWrData;
  wire  sbRamWrEn;
  wire  sbRamRdEn;
  wire [63:0] sbRomRdData;
  wire  dbRdEn;
  wire  dbWrEn;
  wire [33:0] dbRdData;
  reg  dbStateReg;
  reg [31:0] GEN_112;
  wire [33:0] dbResult_data;
  wire [1:0] dbResult_resp;
  wire [4:0] dbReq_addr;
  wire [33:0] dbReq_data;
  wire [1:0] dbReq_op;
  reg [33:0] dbRespReg_data;
  reg [63:0] GEN_113;
  reg [1:0] dbRespReg_resp;
  reg [31:0] GEN_114;
  wire  rdCondWrFailure;
  wire  dbWrNeeded;
  wire [11:0] sbAddr;
  wire [63:0] sbRdData;
  wire [63:0] sbWrData;
  wire [63:0] sbWrMask;
  wire  sbWrEn;
  wire  sbRdEn;
  wire  stallFromDb;
  wire  stallFromSb;
  wire  T_720;
  wire  T_721;
  wire  GEN_11;
  wire  GEN_12;
  wire  T_723;
  wire  T_724;
  wire  T_726;
  wire  T_727;
  wire  GEN_13;
  wire  GEN_14;
  wire  T_731;
  wire  T_732;
  wire  T_733;
  wire  T_735;
  wire  GEN_15;
  wire  GEN_16;
  wire  T_738;
  wire  GEN_17;
  wire  GEN_18;
  wire  T_741;
  wire  T_742;
  wire  T_745;
  wire  GEN_19;
  wire  GEN_20;
  wire  T_750;
  wire  T_751;
  wire  T_754;
  wire  GEN_21;
  wire  GEN_22;
  wire [3:0] T_782;
  wire [2:0] T_783;
  wire [31:0] T_799_0;
  wire [31:0] T_799_1;
  wire [31:0] dbRamWrMask_0;
  wire [31:0] dbRamWrMask_1;
  wire  T_804;
  wire [31:0] T_805;
  wire [31:0] T_806;
  wire [31:0] T_812_0;
  wire [31:0] T_812_1;
  wire [31:0] T_821_0;
  wire [31:0] T_821_1;
  wire [31:0] GEN_0;
  wire [31:0] GEN_23;
  wire [31:0] GEN_24;
  wire [31:0] GEN_1;
  wire [31:0] GEN_25;
  wire [63:0] T_828;
  wire [63:0] T_829;
  wire  T_830;
  wire  T_831;
  wire  T_832;
  wire  T_834;
  wire  T_835;
  wire  T_837;
  wire [63:0] dbRamWrDataVec;
  wire [63:0] T_838;
  wire [63:0] T_839;
  wire [63:0] T_840;
  wire [63:0] T_841;
  wire [63:0] T_842;
  wire [63:0] T_845;
  wire [63:0] T_846;
  wire  T_847;
  wire [2:0] T_848;
  wire [2:0] T_849;
  wire  T_852;
  wire  T_875_interrupt;
  wire  T_875_haltnot;
  wire [9:0] T_875_reserved0;
  wire [2:0] T_875_buserror;
  wire [2:0] T_875_serial;
  wire  T_875_autoincrement;
  wire [2:0] T_875_access;
  wire [9:0] T_875_hartid;
  wire  T_875_ndreset;
  wire  T_875_fullreset;
  wire  T_886;
  wire  T_887;
  wire [9:0] T_888;
  wire [2:0] T_889;
  wire  T_890;
  wire [2:0] T_891;
  wire [2:0] T_892;
  wire [9:0] T_893;
  wire  T_894;
  wire  T_895;
  wire  T_904_interrupt;
  wire  T_904_haltnot;
  wire [31:0] T_904_data;
  wire [31:0] T_908;
  wire  T_913;
  wire  T_915;
  wire  GEN_31;
  wire  T_917;
  wire  T_919;
  wire  T_920;
  wire  GEN_32;
  wire  T_924;
  wire  T_925;
  wire  GEN_33;
  wire  GEN_34;
  wire [9:0] GEN_35;
  wire [2:0] GEN_36;
  wire [2:0] GEN_37;
  wire  GEN_38;
  wire [2:0] GEN_39;
  wire [9:0] GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  T_928;
  wire  T_929;
  wire  T_930;
  wire  GEN_44;
  wire  T_933;
  wire  T_935;
  wire [1:0] T_938;
  wire  T_939;
  wire  T_940;
  wire  GEN_45;
  wire [9:0] GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  T_945;
  wire  GEN_49;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  T_958;
  wire [31:0] GEN_50;
  wire [1:0] T_963;
  wire [33:0] T_964;
  wire [33:0] GEN_51;
  wire [1:0] T_970;
  wire [3:0] T_971;
  wire [13:0] T_972;
  wire [15:0] T_973;
  wire [5:0] T_974;
  wire [1:0] T_975;
  wire [11:0] T_976;
  wire [17:0] T_977;
  wire [33:0] T_978;
  wire [33:0] GEN_53;
  wire  T_980;
  wire  T_986;
  wire [2:0] T_987;
  wire [4:0] T_988;
  wire [3:0] T_989;
  wire [6:0] T_990;
  wire [10:0] T_991;
  wire [15:0] T_992;
  wire [1:0] T_993;
  wire [1:0] T_994;
  wire [3:0] T_995;
  wire [4:0] T_996;
  wire [8:0] T_997;
  wire [13:0] T_998;
  wire [17:0] T_999;
  wire [33:0] T_1000;
  wire [33:0] GEN_54;
  wire  T_1002;
  wire  T_1009;
  wire  T_1010;
  wire  T_1011;
  wire [33:0] GEN_55;
  wire [2:0] T_1013;
  wire  T_1015;
  wire  T_1025;
  wire  T_1026;
  wire  T_1027;
  wire [33:0] GEN_56;
  wire  T_1040;
  wire  T_1041;
  wire [33:0] GEN_57;
  wire  T_1043;
  wire  T_1045;
  wire  T_1046;
  wire  T_1048;
  wire  T_1051;
  wire  T_1052;
  wire  T_1053;
  wire [1:0] T_1056;
  wire  T_1058;
  wire  T_1059;
  wire  T_1061;
  wire  T_1062;
  wire  T_1063;
  wire  T_1064;
  wire  T_1066;
  wire  T_1068;
  wire  GEN_58;
  wire [33:0] GEN_59;
  wire [1:0] GEN_60;
  wire  GEN_61;
  wire [33:0] GEN_62;
  wire [1:0] GEN_63;
  wire  T_1073;
  wire  T_1074;
  wire  GEN_64;
  wire [33:0] GEN_65;
  wire [1:0] GEN_66;
  wire  T_1078;
  wire  T_1079;
  wire  GEN_67;
  wire  GEN_68;
  wire [33:0] GEN_69;
  wire [1:0] GEN_70;
  wire [63:0] T_1101_0;
  wire [63:0] T_1101_1;
  wire [63:0] T_1101_2;
  wire [63:0] T_1101_3;
  wire [63:0] T_1101_4;
  wire [63:0] T_1101_5;
  wire [63:0] T_1101_6;
  wire [63:0] T_1101_7;
  wire [63:0] T_1101_8;
  wire [63:0] T_1101_9;
  wire [63:0] T_1101_10;
  wire [63:0] T_1101_11;
  wire [63:0] T_1101_12;
  wire [63:0] T_1101_13;
  wire [63:0] T_1101_14;
  wire [3:0] T_1104;
  wire [3:0] T_1105;
  wire [63:0] GEN_6;
  wire [63:0] GEN_71;
  wire [63:0] GEN_72;
  wire [63:0] GEN_73;
  wire [63:0] GEN_74;
  wire [63:0] GEN_75;
  wire [63:0] GEN_76;
  wire [63:0] GEN_77;
  wire [63:0] GEN_78;
  wire [63:0] GEN_79;
  wire [63:0] GEN_80;
  wire [63:0] GEN_81;
  wire [63:0] GEN_82;
  wire [63:0] GEN_83;
  wire [63:0] GEN_84;
  wire [31:0] T_1109;
  wire [31:0] T_1110;
  wire [31:0] T_1116_0;
  wire [31:0] T_1116_1;
  wire [31:0] T_1118;
  wire [31:0] T_1119;
  wire [31:0] T_1125_0;
  wire [31:0] T_1125_1;
  wire [31:0] GEN_7;
  wire [31:0] GEN_8;
  wire [3:0] T_1131;
  wire  T_1133;
  wire  GEN_87;
  wire [8:0] T_1134;
  wire  T_1137;
  wire [31:0] GEN_9;
  wire  T_1141;
  wire  T_1142;
  wire  T_1143;
  wire  T_1147;
  wire [31:0] GEN_10;
  wire  T_1151;
  wire  T_1152;
  wire  T_1153;
  wire [63:0] GEN_91;
  wire  GEN_92;
  wire  T_1163;
  wire  T_1164;
  wire  T_1165;
  wire  T_1167;
  wire  T_1168;
  wire [63:0] GEN_93;
  wire  T_1172;
  wire  T_1173;
  wire [63:0] GEN_94;
  reg [25:0] sbAcqReg_addr_block;
  reg [31:0] GEN_115;
  reg [1:0] sbAcqReg_client_xact_id;
  reg [31:0] GEN_116;
  reg [2:0] sbAcqReg_addr_beat;
  reg [31:0] GEN_117;
  reg  sbAcqReg_is_builtin_type;
  reg [31:0] GEN_118;
  reg [2:0] sbAcqReg_a_type;
  reg [31:0] GEN_119;
  reg [10:0] sbAcqReg_union;
  reg [31:0] GEN_120;
  reg [63:0] sbAcqReg_data;
  reg [63:0] GEN_121;
  reg  sbAcqValidReg;
  reg [31:0] GEN_122;
  wire  T_1202;
  wire  sbReg_get;
  wire  T_1203;
  wire  sbReg_getblk;
  wire  T_1204;
  wire  sbReg_put;
  wire  T_1205;
  wire  sbReg_putblk;
  wire  sbMultibeat;
  wire [3:0] T_1207;
  wire [2:0] sbBeatInc1;
  wire  sbLast;
  wire [2:0] T_1216_0;
  wire [2:0] T_1216_1;
  wire  T_1218;
  wire  T_1219;
  wire  T_1220;
  wire  T_1221;
  wire [2:0] T_1222;
  wire [2:0] T_1224;
  wire [28:0] T_1225;
  wire [31:0] T_1226;
  wire  T_1227;
  wire  T_1228;
  wire  T_1229;
  wire  T_1230;
  wire  T_1232;
  wire  T_1233;
  wire  T_1257;
  wire [7:0] T_1258;
  wire [7:0] T_1260;
  wire [7:0] T_1261;
  wire  T_1262;
  wire  T_1263;
  wire  T_1264;
  wire  T_1265;
  wire  T_1266;
  wire  T_1267;
  wire  T_1268;
  wire  T_1269;
  wire [7:0] T_1273;
  wire [7:0] T_1277;
  wire [7:0] T_1281;
  wire [7:0] T_1285;
  wire [7:0] T_1289;
  wire [7:0] T_1293;
  wire [7:0] T_1297;
  wire [7:0] T_1301;
  wire [15:0] T_1302;
  wire [15:0] T_1303;
  wire [31:0] T_1304;
  wire [15:0] T_1305;
  wire [15:0] T_1306;
  wire [31:0] T_1307;
  wire [63:0] T_1308;
  wire  T_1309;
  wire [25:0] GEN_95;
  wire [1:0] GEN_96;
  wire [2:0] GEN_97;
  wire  GEN_98;
  wire [2:0] GEN_99;
  wire [10:0] GEN_100;
  wire [63:0] GEN_101;
  wire  GEN_102;
  wire  T_1311;
  wire  T_1313;
  wire  T_1314;
  wire  GEN_103;
  wire [2:0] GEN_104;
  wire  GEN_105;
  wire  T_1317;
  wire  GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire  T_1335;
  wire [2:0] T_1336;
  wire  T_1337;
  wire [2:0] T_1338;
  wire  T_1339;
  wire [2:0] T_1340;
  wire  T_1341;
  wire [2:0] T_1342;
  wire  T_1343;
  wire [2:0] T_1344;
  wire  T_1345;
  wire [2:0] T_1346;
  wire  T_1347;
  wire [2:0] T_1348;
  wire [2:0] T_1372_addr_beat;
  wire [1:0] T_1372_client_xact_id;
  wire  T_1372_manager_xact_id;
  wire  T_1372_is_builtin_type;
  wire [3:0] T_1372_g_type;
  wire [63:0] T_1372_data;
  wire  T_1397;
  wire  T_1398;
  wire  T_1400;
  wire  T_1401;
  wire  T_1402;
  wire  sbStall;
  wire  T_1404;
  assign io_db_req_ready = T_1064;
  assign io_db_resp_valid = dbStateReg;
  assign io_db_resp_bits_data = dbRespReg_data;
  assign io_db_resp_bits_resp = dbRespReg_resp;
  assign io_debugInterrupts_0 = interruptRegs_0;
  assign io_tl_acquire_ready = T_1404;
  assign io_tl_grant_valid = sbAcqValidReg;
  assign io_tl_grant_bits_addr_beat = T_1372_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_1372_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_1372_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_1372_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_1372_g_type;
  assign io_tl_grant_bits_data = T_1372_data;
  assign io_ndreset = ndresetCtrReg;
  assign io_fullreset = CONTROLReg_fullreset;
  assign CONTROLReset_interrupt = 1'h0;
  assign CONTROLReset_haltnot = 1'h0;
  assign CONTROLReset_reserved0 = 10'h0;
  assign CONTROLReset_buserror = 3'h0;
  assign CONTROLReset_serial = 3'h0;
  assign CONTROLReset_autoincrement = 1'h0;
  assign CONTROLReset_access = 3'h2;
  assign CONTROLReset_hartid = 10'h0;
  assign CONTROLReset_ndreset = 1'h0;
  assign CONTROLReset_fullreset = 1'h0;
  assign CONTROLWrEn = GEN_32;
  assign CONTROLWrData_interrupt = T_875_interrupt;
  assign CONTROLWrData_haltnot = T_875_haltnot;
  assign CONTROLWrData_reserved0 = T_875_reserved0;
  assign CONTROLWrData_buserror = T_875_buserror;
  assign CONTROLWrData_serial = T_875_serial;
  assign CONTROLWrData_autoincrement = T_875_autoincrement;
  assign CONTROLWrData_access = T_875_access;
  assign CONTROLWrData_hartid = T_875_hartid;
  assign CONTROLWrData_ndreset = T_875_ndreset;
  assign CONTROLWrData_fullreset = T_875_fullreset;
  assign CONTROLRdData_interrupt = GEN_2;
  assign CONTROLRdData_haltnot = GEN_3;
  assign CONTROLRdData_reserved0 = CONTROLReg_reserved0;
  assign CONTROLRdData_buserror = CONTROLReg_buserror;
  assign CONTROLRdData_serial = CONTROLReg_serial;
  assign CONTROLRdData_autoincrement = CONTROLReg_autoincrement;
  assign CONTROLRdData_access = CONTROLReg_access;
  assign CONTROLRdData_hartid = CONTROLReg_hartid;
  assign CONTROLRdData_ndreset = ndresetCtrReg;
  assign CONTROLRdData_fullreset = CONTROLReg_fullreset;
  assign DMINFORdData_reserved0 = 2'h0;
  assign DMINFORdData_abussize = 7'h0;
  assign DMINFORdData_serialcount = 4'h0;
  assign DMINFORdData_access128 = 1'h0;
  assign DMINFORdData_access64 = 1'h0;
  assign DMINFORdData_access32 = 1'h0;
  assign DMINFORdData_access16 = 1'h0;
  assign DMINFORdData_accesss8 = 1'h0;
  assign DMINFORdData_dramsize = 6'hf;
  assign DMINFORdData_haltsum = 1'h0;
  assign DMINFORdData_reserved1 = 3'h0;
  assign DMINFORdData_authenticated = 1'h1;
  assign DMINFORdData_authbusy = 1'h0;
  assign DMINFORdData_authtype = 2'h0;
  assign DMINFORdData_version = 2'h1;
  assign HALTSUMRdData_serialfull = 1'h0;
  assign HALTSUMRdData_serialvalid = 1'h0;
  assign HALTSUMRdData_acks = {{31'd0}, haltnotSummary};
  assign RAMWrData_interrupt = T_904_interrupt;
  assign RAMWrData_haltnot = T_904_haltnot;
  assign RAMWrData_data = T_904_data;
  assign RAMRdData_interrupt = GEN_4;
  assign RAMRdData_haltnot = GEN_5;
  assign RAMRdData_data = dbRamRdData;
  assign SETHALTNOTWrEn = T_1143;
  assign SETHALTNOTWrData = GEN_7[9:0];
  assign CLEARDEBINTWrEn = T_1153;
  assign CLEARDEBINTWrData = GEN_8[9:0];
  assign T_655_0 = 1'h0;
  assign T_666_0 = 1'h0;
  assign haltnotStatus_0 = {{31'd0}, haltnotRegs_0};
  assign rdHaltnotStatus = GEN_50;
  assign haltnotSummary = haltnotStatus_0 != 32'h0;
  assign ramMem_T_850_addr = ramAddr;
  assign ramMem_T_850_en = 1'h1;
  assign ramMem_T_850_data = ramMem[ramMem_T_850_addr];
  assign ramMem_T_851_data = ramWrData;
  assign ramMem_T_851_addr = ramAddr;
  assign ramMem_T_851_mask = ramWrEn;
  assign ramMem_T_851_en = ramWrEn;
  assign ramAddr = T_849;
  assign ramRdData = ramMem_T_850_data;
  assign ramWrData = T_846;
  assign ramWrMask = T_829;
  assign ramWrEn = T_852;
  assign dbRamAddr = T_782;
  assign dbRamRdData = GEN_1;
  assign dbRamWrData = dbReq_data[31:0];
  assign dbRamWrEn = GEN_31;
  assign dbRamRdEn = 1'h0;
  assign sbRamAddr = T_783;
  assign sbRamRdData = ramRdData;
  assign sbRamWrData = sbWrData;
  assign sbRamWrEn = GEN_87;
  assign sbRamRdEn = GEN_92;
  assign sbRomRdData = GEN_6;
  assign dbRdEn = T_1066;
  assign dbWrEn = T_1068;
  assign dbRdData = GEN_57;
  assign dbResult_data = dbRdData;
  assign dbResult_resp = T_1056;
  assign dbReq_addr = io_db_req_bits_addr;
  assign dbReq_data = io_db_req_bits_data;
  assign dbReq_op = io_db_req_bits_op;
  assign rdCondWrFailure = T_1046;
  assign dbWrNeeded = T_1053;
  assign sbAddr = T_1226[11:0];
  assign sbRdData = GEN_94;
  assign sbWrData = sbAcqReg_data;
  assign sbWrMask = T_1308;
  assign sbWrEn = T_1230;
  assign sbRdEn = T_1228;
  assign stallFromDb = 1'h0;
  assign stallFromSb = T_831;
  assign T_720 = CONTROLWrData_hartid == 10'h0;
  assign T_721 = interruptRegs_0 | CONTROLWrData_interrupt;
  assign GEN_11 = T_720 ? T_721 : interruptRegs_0;
  assign GEN_12 = CONTROLWrEn ? GEN_11 : interruptRegs_0;
  assign T_723 = CONTROLWrEn == 1'h0;
  assign T_724 = T_723 & dbRamWrEn;
  assign T_726 = CONTROLReg_hartid == 10'h0;
  assign T_727 = interruptRegs_0 | RAMWrData_interrupt;
  assign GEN_13 = T_726 ? T_727 : GEN_12;
  assign GEN_14 = T_724 ? GEN_13 : GEN_12;
  assign T_731 = dbRamWrEn == 1'h0;
  assign T_732 = T_723 & T_731;
  assign T_733 = T_732 & CLEARDEBINTWrEn;
  assign T_735 = CLEARDEBINTWrData == 10'h0;
  assign GEN_15 = T_735 ? 1'h0 : GEN_14;
  assign GEN_16 = T_733 ? GEN_15 : GEN_14;
  assign T_738 = SETHALTNOTWrData == 10'h0;
  assign GEN_17 = T_738 ? 1'h1 : haltnotRegs_0;
  assign GEN_18 = SETHALTNOTWrEn ? GEN_17 : haltnotRegs_0;
  assign T_741 = SETHALTNOTWrEn == 1'h0;
  assign T_742 = T_741 & CONTROLWrEn;
  assign T_745 = haltnotRegs_0 & CONTROLWrData_haltnot;
  assign GEN_19 = T_720 ? T_745 : GEN_18;
  assign GEN_20 = T_742 ? GEN_19 : GEN_18;
  assign T_750 = T_741 & T_723;
  assign T_751 = T_750 & dbRamWrEn;
  assign T_754 = haltnotRegs_0 & RAMWrData_haltnot;
  assign GEN_21 = T_726 ? T_754 : GEN_20;
  assign GEN_22 = T_751 ? GEN_21 : GEN_20;
  assign T_782 = dbReq_addr[3:0];
  assign T_783 = sbAddr[5:3];
  assign T_799_0 = 32'hffffffff;
  assign T_799_1 = 32'hffffffff;
  assign dbRamWrMask_0 = GEN_23;
  assign dbRamWrMask_1 = GEN_24;
  assign T_804 = dbRamAddr[0];
  assign T_805 = ramRdData[31:0];
  assign T_806 = ramRdData[63:32];
  assign T_812_0 = T_805;
  assign T_812_1 = T_806;
  assign T_821_0 = 32'h0;
  assign T_821_1 = 32'h0;
  assign GEN_0 = 32'hffffffff;
  assign GEN_23 = 1'h0 == T_804 ? GEN_0 : T_821_0;
  assign GEN_24 = T_804 ? GEN_0 : T_821_1;
  assign GEN_1 = GEN_25;
  assign GEN_25 = T_804 ? T_812_1 : T_812_0;
  assign T_828 = {dbRamWrMask_1,dbRamWrMask_0};
  assign T_829 = sbRamWrEn ? sbWrMask : T_828;
  assign T_830 = dbRamWrEn | dbRamRdEn;
  assign T_831 = sbRamRdEn | sbRamWrEn;
  assign T_832 = T_830 & T_831;
  assign T_834 = T_832 == 1'h0;
  assign T_835 = T_834 | reset;
  assign T_837 = T_835 == 1'h0;
  assign dbRamWrDataVec = {dbRamWrData,dbRamWrData};
  assign T_838 = ramWrMask & sbRamWrData;
  assign T_839 = ~ ramWrMask;
  assign T_840 = T_839 & ramRdData;
  assign T_841 = T_838 | T_840;
  assign T_842 = ramWrMask & dbRamWrDataVec;
  assign T_845 = T_842 | T_840;
  assign T_846 = sbRamWrEn ? T_841 : T_845;
  assign T_847 = sbRamWrEn | sbRamRdEn;
  assign T_848 = dbRamAddr[3:1];
  assign T_849 = T_847 ? sbRamAddr : T_848;
  assign T_852 = sbRamWrEn | dbRamWrEn;
  assign T_875_interrupt = T_895;
  assign T_875_haltnot = T_894;
  assign T_875_reserved0 = T_893;
  assign T_875_buserror = T_892;
  assign T_875_serial = T_891;
  assign T_875_autoincrement = T_890;
  assign T_875_access = T_889;
  assign T_875_hartid = T_888;
  assign T_875_ndreset = T_887;
  assign T_875_fullreset = T_886;
  assign T_886 = dbReq_data[0];
  assign T_887 = dbReq_data[1];
  assign T_888 = dbReq_data[11:2];
  assign T_889 = dbReq_data[14:12];
  assign T_890 = dbReq_data[15];
  assign T_891 = dbReq_data[18:16];
  assign T_892 = dbReq_data[21:19];
  assign T_893 = dbReq_data[31:22];
  assign T_894 = dbReq_data[32];
  assign T_895 = dbReq_data[33];
  assign T_904_interrupt = T_895;
  assign T_904_haltnot = T_894;
  assign T_904_data = T_908;
  assign T_908 = dbReq_data[31:0];
  assign T_913 = dbReq_addr[4:4];
  assign T_915 = T_913 == 1'h0;
  assign GEN_31 = T_915 ? dbWrEn : 1'h0;
  assign T_917 = dbReq_addr == 5'h10;
  assign T_919 = T_915 == 1'h0;
  assign T_920 = T_919 & T_917;
  assign GEN_32 = T_920 ? dbWrEn : 1'h0;
  assign T_924 = T_917 == 1'h0;
  assign T_925 = T_919 & T_924;
  assign GEN_33 = reset ? CONTROLReset_interrupt : CONTROLReg_interrupt;
  assign GEN_34 = reset ? CONTROLReset_haltnot : CONTROLReg_haltnot;
  assign GEN_35 = reset ? CONTROLReset_reserved0 : CONTROLReg_reserved0;
  assign GEN_36 = reset ? CONTROLReset_buserror : CONTROLReg_buserror;
  assign GEN_37 = reset ? CONTROLReset_serial : CONTROLReg_serial;
  assign GEN_38 = reset ? CONTROLReset_autoincrement : CONTROLReg_autoincrement;
  assign GEN_39 = reset ? CONTROLReset_access : CONTROLReg_access;
  assign GEN_40 = reset ? CONTROLReset_hartid : CONTROLReg_hartid;
  assign GEN_41 = reset ? CONTROLReset_ndreset : CONTROLReg_ndreset;
  assign GEN_42 = reset ? CONTROLReset_fullreset : CONTROLReg_fullreset;
  assign GEN_43 = reset ? 1'h0 : ndresetCtrReg;
  assign T_928 = reset == 1'h0;
  assign T_929 = T_928 & CONTROLWrEn;
  assign T_930 = CONTROLReg_fullreset | CONTROLWrData_fullreset;
  assign GEN_44 = CONTROLWrData_ndreset ? 1'h1 : GEN_43;
  assign T_933 = CONTROLWrData_ndreset == 1'h0;
  assign T_935 = ndresetCtrReg == 1'h0;
  assign T_938 = ndresetCtrReg - 1'h1;
  assign T_939 = T_938[0:0];
  assign T_940 = T_935 ? 1'h0 : T_939;
  assign GEN_45 = T_933 ? T_940 : GEN_44;
  assign GEN_46 = T_929 ? CONTROLWrData_hartid : GEN_40;
  assign GEN_47 = T_929 ? T_930 : GEN_42;
  assign GEN_48 = T_929 ? GEN_45 : GEN_43;
  assign T_945 = T_928 & T_723;
  assign GEN_49 = T_945 ? T_940 : GEN_48;
  assign GEN_2 = interruptRegs_0;
  assign GEN_3 = haltnotRegs_0;
  assign GEN_4 = interruptRegs_0;
  assign GEN_5 = haltnotRegs_0;
  assign T_958 = dbReq_addr == 5'h0;
  assign GEN_50 = T_958 ? haltnotStatus_0 : 32'h0;
  assign T_963 = {RAMRdData_interrupt,RAMRdData_haltnot};
  assign T_964 = {T_963,RAMRdData_data};
  assign GEN_51 = T_915 ? T_964 : 34'h0;
  assign T_970 = {CONTROLRdData_ndreset,CONTROLRdData_fullreset};
  assign T_971 = {CONTROLRdData_autoincrement,CONTROLRdData_access};
  assign T_972 = {T_971,CONTROLRdData_hartid};
  assign T_973 = {T_972,T_970};
  assign T_974 = {CONTROLRdData_buserror,CONTROLRdData_serial};
  assign T_975 = {CONTROLRdData_interrupt,CONTROLRdData_haltnot};
  assign T_976 = {T_975,CONTROLRdData_reserved0};
  assign T_977 = {T_976,T_974};
  assign T_978 = {T_977,T_973};
  assign GEN_53 = T_920 ? T_978 : GEN_51;
  assign T_980 = dbReq_addr == 5'h11;
  assign T_986 = T_925 & T_980;
  assign T_987 = {DMINFORdData_authbusy,DMINFORdData_authtype};
  assign T_988 = {T_987,DMINFORdData_version};
  assign T_989 = {DMINFORdData_reserved1,DMINFORdData_authenticated};
  assign T_990 = {DMINFORdData_dramsize,DMINFORdData_haltsum};
  assign T_991 = {T_990,T_989};
  assign T_992 = {T_991,T_988};
  assign T_993 = {DMINFORdData_access16,DMINFORdData_accesss8};
  assign T_994 = {DMINFORdData_access64,DMINFORdData_access32};
  assign T_995 = {T_994,T_993};
  assign T_996 = {DMINFORdData_serialcount,DMINFORdData_access128};
  assign T_997 = {DMINFORdData_reserved0,DMINFORdData_abussize};
  assign T_998 = {T_997,T_996};
  assign T_999 = {T_998,T_995};
  assign T_1000 = {T_999,T_992};
  assign GEN_54 = T_986 ? T_1000 : GEN_53;
  assign T_1002 = dbReq_addr == 5'h1b;
  assign T_1009 = T_980 == 1'h0;
  assign T_1010 = T_925 & T_1009;
  assign T_1011 = T_1010 & T_1002;
  assign GEN_55 = T_1011 ? 34'h0 : GEN_54;
  assign T_1013 = dbReq_addr[4:2];
  assign T_1015 = T_1013 == 3'h7;
  assign T_1025 = T_1002 == 1'h0;
  assign T_1026 = T_1010 & T_1025;
  assign T_1027 = T_1026 & T_1015;
  assign GEN_56 = T_1027 ? {{2'd0}, rdHaltnotStatus} : GEN_55;
  assign T_1040 = T_1015 == 1'h0;
  assign T_1041 = T_1026 & T_1040;
  assign GEN_57 = T_1041 ? 34'h0 : GEN_56;
  assign T_1043 = dbRdData[33];
  assign T_1045 = dbReq_op == 2'h3;
  assign T_1046 = T_1043 & T_1045;
  assign T_1048 = dbReq_op == 2'h2;
  assign T_1051 = ~ rdCondWrFailure;
  assign T_1052 = T_1045 & T_1051;
  assign T_1053 = T_1048 | T_1052;
  assign T_1056 = rdCondWrFailure ? 2'h1 : 2'h0;
  assign T_1058 = stallFromSb == 1'h0;
  assign T_1059 = dbStateReg == 1'h0;
  assign T_1061 = io_db_resp_ready & io_db_resp_valid;
  assign T_1062 = dbStateReg & T_1061;
  assign T_1063 = T_1059 | T_1062;
  assign T_1064 = T_1058 & T_1063;
  assign T_1066 = io_db_req_ready & io_db_req_valid;
  assign T_1068 = dbWrNeeded & T_1066;
  assign GEN_58 = T_1066 ? 1'h1 : dbStateReg;
  assign GEN_59 = T_1066 ? dbResult_data : dbRespReg_data;
  assign GEN_60 = T_1066 ? dbResult_resp : dbRespReg_resp;
  assign GEN_61 = T_1059 ? GEN_58 : dbStateReg;
  assign GEN_62 = T_1059 ? GEN_59 : dbRespReg_data;
  assign GEN_63 = T_1059 ? GEN_60 : dbRespReg_resp;
  assign T_1073 = T_1059 == 1'h0;
  assign T_1074 = T_1073 & dbStateReg;
  assign GEN_64 = T_1066 ? 1'h1 : GEN_61;
  assign GEN_65 = T_1066 ? dbResult_data : GEN_62;
  assign GEN_66 = T_1066 ? dbResult_resp : GEN_63;
  assign T_1078 = T_1066 == 1'h0;
  assign T_1079 = T_1078 & T_1061;
  assign GEN_67 = T_1079 ? 1'h0 : GEN_64;
  assign GEN_68 = T_1074 ? GEN_67 : GEN_61;
  assign GEN_69 = T_1074 ? GEN_65 : GEN_62;
  assign GEN_70 = T_1074 ? GEN_66 : GEN_63;
  assign T_1101_0 = 64'hc0006f03c0006f;
  assign T_1101_1 = 64'h80006ffff00413;
  assign T_1101_2 = 64'hff0000f00000413;
  assign T_1101_3 = 64'h42802e2343803483;
  assign T_1101_4 = 64'h10802023f1402473;
  assign T_1101_5 = 64'h8474137b002473;
  assign T_1101_6 = 64'h7b20247302041a63;
  assign T_1101_7 = 64'h7b2410737b200073;
  assign T_1101_8 = 64'h1c0474137b002473;
  assign T_1101_9 = 64'h41663f4040413;
  assign T_1101_10 = 64'h4000006742903c23;
  assign T_1101_11 = 64'h10802623f1402473;
  assign T_1101_12 = 64'h7b0024737b046073;
  assign T_1101_13 = 64'hfe040ce302047413;
  assign T_1101_14 = 64'hfe1ff06f;
  assign T_1104 = T_1105;
  assign T_1105 = sbAddr[6:3];
  assign GEN_6 = GEN_84;
  assign GEN_71 = 4'h1 == T_1104 ? T_1101_1 : T_1101_0;
  assign GEN_72 = 4'h2 == T_1104 ? T_1101_2 : GEN_71;
  assign GEN_73 = 4'h3 == T_1104 ? T_1101_3 : GEN_72;
  assign GEN_74 = 4'h4 == T_1104 ? T_1101_4 : GEN_73;
  assign GEN_75 = 4'h5 == T_1104 ? T_1101_5 : GEN_74;
  assign GEN_76 = 4'h6 == T_1104 ? T_1101_6 : GEN_75;
  assign GEN_77 = 4'h7 == T_1104 ? T_1101_7 : GEN_76;
  assign GEN_78 = 4'h8 == T_1104 ? T_1101_8 : GEN_77;
  assign GEN_79 = 4'h9 == T_1104 ? T_1101_9 : GEN_78;
  assign GEN_80 = 4'ha == T_1104 ? T_1101_10 : GEN_79;
  assign GEN_81 = 4'hb == T_1104 ? T_1101_11 : GEN_80;
  assign GEN_82 = 4'hc == T_1104 ? T_1101_12 : GEN_81;
  assign GEN_83 = 4'hd == T_1104 ? T_1101_13 : GEN_82;
  assign GEN_84 = 4'he == T_1104 ? T_1101_14 : GEN_83;
  assign T_1109 = sbWrData[31:0];
  assign T_1110 = sbWrData[63:32];
  assign T_1116_0 = T_1109;
  assign T_1116_1 = T_1110;
  assign T_1118 = sbWrMask[31:0];
  assign T_1119 = sbWrMask[63:32];
  assign T_1125_0 = T_1118;
  assign T_1125_1 = T_1119;
  assign GEN_7 = T_1116_1;
  assign GEN_8 = T_1116_0;
  assign T_1131 = sbAddr[11:8];
  assign T_1133 = T_1131 == 4'h4;
  assign GEN_87 = T_1133 ? sbWrEn : 1'h0;
  assign T_1134 = sbAddr[11:3];
  assign T_1137 = T_1134 == 9'h21;
  assign GEN_9 = T_1125_1;
  assign T_1141 = GEN_9 != 32'h0;
  assign T_1142 = T_1137 & T_1141;
  assign T_1143 = T_1142 & sbWrEn;
  assign T_1147 = T_1134 == 9'h20;
  assign GEN_10 = T_1125_0;
  assign T_1151 = GEN_10 != 32'h0;
  assign T_1152 = T_1147 & T_1151;
  assign T_1153 = T_1152 & sbWrEn;
  assign GEN_91 = T_1133 ? sbRamRdData : 64'h0;
  assign GEN_92 = T_1133 ? sbRdEn : 1'h0;
  assign T_1163 = T_1131 == 4'h8;
  assign T_1164 = T_1131 == 4'h9;
  assign T_1165 = T_1163 | T_1164;
  assign T_1167 = T_1133 == 1'h0;
  assign T_1168 = T_1167 & T_1165;
  assign GEN_93 = T_1168 ? sbRomRdData : GEN_91;
  assign T_1172 = T_1165 == 1'h0;
  assign T_1173 = T_1167 & T_1172;
  assign GEN_94 = T_1173 ? 64'h0 : GEN_93;
  assign T_1202 = sbAcqReg_a_type == 3'h0;
  assign sbReg_get = sbAcqReg_is_builtin_type & T_1202;
  assign T_1203 = sbAcqReg_a_type == 3'h1;
  assign sbReg_getblk = sbAcqReg_is_builtin_type & T_1203;
  assign T_1204 = sbAcqReg_a_type == 3'h2;
  assign sbReg_put = sbAcqReg_is_builtin_type & T_1204;
  assign T_1205 = sbAcqReg_a_type == 3'h3;
  assign sbReg_putblk = sbAcqReg_is_builtin_type & T_1205;
  assign sbMultibeat = sbReg_getblk & sbAcqValidReg;
  assign T_1207 = sbAcqReg_addr_beat + 3'h1;
  assign sbBeatInc1 = T_1207[2:0];
  assign sbLast = sbAcqReg_addr_beat == 3'h7;
  assign T_1216_0 = 3'h0;
  assign T_1216_1 = 3'h4;
  assign T_1218 = sbAcqReg_a_type == T_1216_0;
  assign T_1219 = sbAcqReg_a_type == T_1216_1;
  assign T_1220 = T_1218 | T_1219;
  assign T_1221 = sbAcqReg_is_builtin_type & T_1220;
  assign T_1222 = sbAcqReg_union[10:8];
  assign T_1224 = T_1221 ? T_1222 : 3'h0;
  assign T_1225 = {sbAcqReg_addr_block,sbAcqReg_addr_beat};
  assign T_1226 = {T_1225,T_1224};
  assign T_1227 = sbReg_get | sbReg_getblk;
  assign T_1228 = sbAcqValidReg & T_1227;
  assign T_1229 = sbReg_put | sbReg_putblk;
  assign T_1230 = sbAcqValidReg & T_1229;
  assign T_1232 = sbAcqReg_a_type == 3'h4;
  assign T_1233 = sbAcqReg_is_builtin_type & T_1232;
  assign T_1257 = sbReg_putblk | sbReg_put;
  assign T_1258 = sbAcqReg_union[8:1];
  assign T_1260 = T_1257 ? T_1258 : 8'h0;
  assign T_1261 = T_1233 ? 8'hff : T_1260;
  assign T_1262 = T_1261[0];
  assign T_1263 = T_1261[1];
  assign T_1264 = T_1261[2];
  assign T_1265 = T_1261[3];
  assign T_1266 = T_1261[4];
  assign T_1267 = T_1261[5];
  assign T_1268 = T_1261[6];
  assign T_1269 = T_1261[7];
  assign T_1273 = T_1262 ? 8'hff : 8'h0;
  assign T_1277 = T_1263 ? 8'hff : 8'h0;
  assign T_1281 = T_1264 ? 8'hff : 8'h0;
  assign T_1285 = T_1265 ? 8'hff : 8'h0;
  assign T_1289 = T_1266 ? 8'hff : 8'h0;
  assign T_1293 = T_1267 ? 8'hff : 8'h0;
  assign T_1297 = T_1268 ? 8'hff : 8'h0;
  assign T_1301 = T_1269 ? 8'hff : 8'h0;
  assign T_1302 = {T_1277,T_1273};
  assign T_1303 = {T_1285,T_1281};
  assign T_1304 = {T_1303,T_1302};
  assign T_1305 = {T_1293,T_1289};
  assign T_1306 = {T_1301,T_1297};
  assign T_1307 = {T_1306,T_1305};
  assign T_1308 = {T_1307,T_1304};
  assign T_1309 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign GEN_95 = T_1309 ? io_tl_acquire_bits_addr_block : sbAcqReg_addr_block;
  assign GEN_96 = T_1309 ? io_tl_acquire_bits_client_xact_id : sbAcqReg_client_xact_id;
  assign GEN_97 = T_1309 ? io_tl_acquire_bits_addr_beat : sbAcqReg_addr_beat;
  assign GEN_98 = T_1309 ? io_tl_acquire_bits_is_builtin_type : sbAcqReg_is_builtin_type;
  assign GEN_99 = T_1309 ? io_tl_acquire_bits_a_type : sbAcqReg_a_type;
  assign GEN_100 = T_1309 ? io_tl_acquire_bits_union : sbAcqReg_union;
  assign GEN_101 = T_1309 ? io_tl_acquire_bits_data : sbAcqReg_data;
  assign GEN_102 = T_1309 ? 1'h1 : sbAcqValidReg;
  assign T_1311 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_1313 = T_1309 == 1'h0;
  assign T_1314 = T_1313 & T_1311;
  assign GEN_103 = sbLast ? 1'h0 : GEN_102;
  assign GEN_104 = sbMultibeat ? sbBeatInc1 : GEN_97;
  assign GEN_105 = sbMultibeat ? GEN_103 : GEN_102;
  assign T_1317 = sbMultibeat == 1'h0;
  assign GEN_106 = T_1317 ? 1'h0 : GEN_105;
  assign GEN_107 = T_1314 ? GEN_104 : GEN_97;
  assign GEN_108 = T_1314 ? GEN_106 : GEN_102;
  assign T_1335 = 3'h6 == sbAcqReg_a_type;
  assign T_1336 = T_1335 ? 3'h1 : 3'h3;
  assign T_1337 = 3'h5 == sbAcqReg_a_type;
  assign T_1338 = T_1337 ? 3'h1 : T_1336;
  assign T_1339 = 3'h4 == sbAcqReg_a_type;
  assign T_1340 = T_1339 ? 3'h4 : T_1338;
  assign T_1341 = 3'h3 == sbAcqReg_a_type;
  assign T_1342 = T_1341 ? 3'h3 : T_1340;
  assign T_1343 = 3'h2 == sbAcqReg_a_type;
  assign T_1344 = T_1343 ? 3'h3 : T_1342;
  assign T_1345 = 3'h1 == sbAcqReg_a_type;
  assign T_1346 = T_1345 ? 3'h5 : T_1344;
  assign T_1347 = 3'h0 == sbAcqReg_a_type;
  assign T_1348 = T_1347 ? 3'h4 : T_1346;
  assign T_1372_addr_beat = sbAcqReg_addr_beat;
  assign T_1372_client_xact_id = sbAcqReg_client_xact_id;
  assign T_1372_manager_xact_id = 1'h0;
  assign T_1372_is_builtin_type = 1'h1;
  assign T_1372_g_type = {{1'd0}, T_1348};
  assign T_1372_data = sbRdData;
  assign T_1397 = sbLast == 1'h0;
  assign T_1398 = sbMultibeat & T_1397;
  assign T_1400 = io_tl_grant_ready == 1'h0;
  assign T_1401 = io_tl_grant_valid & T_1400;
  assign T_1402 = T_1398 | T_1401;
  assign sbStall = T_1402 | stallFromDb;
  assign T_1404 = sbStall == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_26 = {1{$random}};
  CONTROLReg_interrupt = GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_27 = {1{$random}};
  CONTROLReg_haltnot = GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_28 = {1{$random}};
  CONTROLReg_reserved0 = GEN_28[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  CONTROLReg_buserror = GEN_29[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  CONTROLReg_serial = GEN_30[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  CONTROLReg_autoincrement = GEN_52[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {1{$random}};
  CONTROLReg_access = GEN_85[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  CONTROLReg_hartid = GEN_86[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  CONTROLReg_ndreset = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {1{$random}};
  CONTROLReg_fullreset = GEN_89[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {1{$random}};
  ndresetCtrReg = GEN_90[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_109 = {1{$random}};
  interruptRegs_0 = GEN_109[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_110 = {1{$random}};
  haltnotRegs_0 = GEN_110[0:0];
  `endif
  GEN_111 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ramMem[initvar] = GEN_111[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {1{$random}};
  dbStateReg = GEN_112[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_113 = {2{$random}};
  dbRespReg_data = GEN_113[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_114 = {1{$random}};
  dbRespReg_resp = GEN_114[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  sbAcqReg_addr_block = GEN_115[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_116 = {1{$random}};
  sbAcqReg_client_xact_id = GEN_116[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_117 = {1{$random}};
  sbAcqReg_addr_beat = GEN_117[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_118 = {1{$random}};
  sbAcqReg_is_builtin_type = GEN_118[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  sbAcqReg_a_type = GEN_119[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  sbAcqReg_union = GEN_120[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_121 = {2{$random}};
  sbAcqReg_data = GEN_121[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_122 = {1{$random}};
  sbAcqValidReg = GEN_122[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_interrupt <= CONTROLReset_interrupt;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_haltnot <= CONTROLReset_haltnot;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_reserved0 <= CONTROLReset_reserved0;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_buserror <= CONTROLReset_buserror;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_serial <= CONTROLReset_serial;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_autoincrement <= CONTROLReset_autoincrement;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_access <= CONTROLReset_access;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_929) begin
        CONTROLReg_hartid <= CONTROLWrData_hartid;
      end else begin
        if(reset) begin
          CONTROLReg_hartid <= CONTROLReset_hartid;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_ndreset <= CONTROLReset_ndreset;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_929) begin
        CONTROLReg_fullreset <= T_930;
      end else begin
        if(reset) begin
          CONTROLReg_fullreset <= CONTROLReset_fullreset;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_945) begin
        if(T_935) begin
          ndresetCtrReg <= 1'h0;
        end else begin
          ndresetCtrReg <= T_939;
        end
      end else begin
        if(T_929) begin
          if(T_933) begin
            if(T_935) begin
              ndresetCtrReg <= 1'h0;
            end else begin
              ndresetCtrReg <= T_939;
            end
          end else begin
            if(CONTROLWrData_ndreset) begin
              ndresetCtrReg <= 1'h1;
            end else begin
              if(reset) begin
                ndresetCtrReg <= 1'h0;
              end
            end
          end
        end else begin
          if(reset) begin
            ndresetCtrReg <= 1'h0;
          end
        end
      end
    end
    if(reset) begin
      interruptRegs_0 <= T_655_0;
    end else begin
      if(T_733) begin
        if(T_735) begin
          interruptRegs_0 <= 1'h0;
        end else begin
          if(T_724) begin
            if(T_726) begin
              interruptRegs_0 <= T_727;
            end else begin
              if(CONTROLWrEn) begin
                if(T_720) begin
                  interruptRegs_0 <= T_721;
                end
              end
            end
          end else begin
            if(CONTROLWrEn) begin
              if(T_720) begin
                interruptRegs_0 <= T_721;
              end
            end
          end
        end
      end else begin
        if(T_724) begin
          if(T_726) begin
            interruptRegs_0 <= T_727;
          end else begin
            if(CONTROLWrEn) begin
              if(T_720) begin
                interruptRegs_0 <= T_721;
              end
            end
          end
        end else begin
          if(CONTROLWrEn) begin
            if(T_720) begin
              interruptRegs_0 <= T_721;
            end
          end
        end
      end
    end
    if(reset) begin
      haltnotRegs_0 <= T_666_0;
    end else begin
      if(T_751) begin
        if(T_726) begin
          haltnotRegs_0 <= T_754;
        end else begin
          if(T_742) begin
            if(T_720) begin
              haltnotRegs_0 <= T_745;
            end else begin
              if(SETHALTNOTWrEn) begin
                if(T_738) begin
                  haltnotRegs_0 <= 1'h1;
                end
              end
            end
          end else begin
            if(SETHALTNOTWrEn) begin
              if(T_738) begin
                haltnotRegs_0 <= 1'h1;
              end
            end
          end
        end
      end else begin
        if(T_742) begin
          if(T_720) begin
            haltnotRegs_0 <= T_745;
          end else begin
            if(SETHALTNOTWrEn) begin
              if(T_738) begin
                haltnotRegs_0 <= 1'h1;
              end
            end
          end
        end else begin
          if(SETHALTNOTWrEn) begin
            if(T_738) begin
              haltnotRegs_0 <= 1'h1;
            end
          end
        end
      end
    end
    if(ramMem_T_851_en & ramMem_T_851_mask) begin
      ramMem[ramMem_T_851_addr] <= ramMem_T_851_data;
    end
    if(reset) begin
      dbStateReg <= 1'h0;
    end else begin
      if(T_1074) begin
        if(T_1079) begin
          dbStateReg <= 1'h0;
        end else begin
          if(T_1066) begin
            dbStateReg <= 1'h1;
          end else begin
            if(T_1059) begin
              if(T_1066) begin
                dbStateReg <= 1'h1;
              end
            end
          end
        end
      end else begin
        if(T_1059) begin
          if(T_1066) begin
            dbStateReg <= 1'h1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1074) begin
        if(T_1066) begin
          dbRespReg_data <= dbResult_data;
        end else begin
          if(T_1059) begin
            if(T_1066) begin
              dbRespReg_data <= dbResult_data;
            end
          end
        end
      end else begin
        if(T_1059) begin
          if(T_1066) begin
            dbRespReg_data <= dbResult_data;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1074) begin
        if(T_1066) begin
          dbRespReg_resp <= dbResult_resp;
        end else begin
          if(T_1059) begin
            if(T_1066) begin
              dbRespReg_resp <= dbResult_resp;
            end
          end
        end
      end else begin
        if(T_1059) begin
          if(T_1066) begin
            dbRespReg_resp <= dbResult_resp;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_addr_block <= io_tl_acquire_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_client_xact_id <= io_tl_acquire_bits_client_xact_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1314) begin
        if(sbMultibeat) begin
          sbAcqReg_addr_beat <= sbBeatInc1;
        end else begin
          if(T_1309) begin
            sbAcqReg_addr_beat <= io_tl_acquire_bits_addr_beat;
          end
        end
      end else begin
        if(T_1309) begin
          sbAcqReg_addr_beat <= io_tl_acquire_bits_addr_beat;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_is_builtin_type <= io_tl_acquire_bits_is_builtin_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_a_type <= io_tl_acquire_bits_a_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_union <= io_tl_acquire_bits_union;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_data <= io_tl_acquire_bits_data;
      end
    end
    if(reset) begin
      sbAcqValidReg <= 1'h0;
    end else begin
      if(T_1314) begin
        if(T_1317) begin
          sbAcqValidReg <= 1'h0;
        end else begin
          if(sbMultibeat) begin
            if(sbLast) begin
              sbAcqValidReg <= 1'h0;
            end else begin
              if(T_1309) begin
                sbAcqValidReg <= 1'h1;
              end
            end
          end else begin
            if(T_1309) begin
              sbAcqValidReg <= 1'h1;
            end
          end
        end
      end else begin
        if(T_1309) begin
          sbAcqValidReg <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_837) begin
          $fwrite(32'h80000002,"Assertion failed: Stall logic should have prevented concurrent SB/DB RAM Access\n    at Debug.scala:650 assert (!((dbRamWrEn | dbRamRdEn) & (sbRamRdEn | sbRamWrEn)), \"Stall logic should have prevented concurrent SB/DB RAM Access\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_837) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module PRCI(
  input   clk,
  input   reset,
  input   io_interrupts_0_meip,
  input   io_interrupts_0_seip,
  input   io_interrupts_0_debug,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [10:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_tiles_0_reset,
  output  io_tiles_0_id,
  output  io_tiles_0_interrupts_meip,
  output  io_tiles_0_interrupts_seip,
  output  io_tiles_0_interrupts_debug,
  output  io_tiles_0_interrupts_mtip,
  output  io_tiles_0_interrupts_msip,
  input   io_rtcTick
);
  reg [63:0] timecmp_0;
  reg [63:0] GEN_3;
  reg [63:0] time$;
  reg [63:0] GEN_4;
  wire [64:0] T_525;
  wire [63:0] T_526;
  wire [63:0] GEN_0;
  wire [31:0] T_533_0;
  reg [31:0] ipi_0;
  reg [31:0] GEN_5;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [10:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [10:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire [2:0] T_568_0;
  wire [2:0] T_568_1;
  wire  T_570;
  wire  T_571;
  wire  T_572;
  wire  T_573;
  wire [2:0] T_574;
  wire [2:0] T_576;
  wire [28:0] T_577;
  wire [31:0] T_578;
  wire [15:0] addr;
  wire [63:0] rdata;
  wire  T_598;
  wire [2:0] T_599;
  wire  T_600;
  wire [2:0] T_601;
  wire  T_602;
  wire [2:0] T_603;
  wire  T_604;
  wire [2:0] T_605;
  wire  T_606;
  wire [2:0] T_607;
  wire  T_608;
  wire [2:0] T_609;
  wire  T_610;
  wire [2:0] T_611;
  wire [2:0] T_636_addr_beat;
  wire [1:0] T_636_client_xact_id;
  wire  T_636_manager_xact_id;
  wire  T_636_is_builtin_type;
  wire [3:0] T_636_g_type;
  wire [63:0] T_636_data;
  wire  T_658;
  wire  T_659;
  wire [2:0] T_667_0;
  wire [2:0] T_667_1;
  wire [2:0] T_685_0;
  wire [2:0] T_685_1;
  wire  T_697;
  wire  T_698;
  wire  T_717;
  wire  T_718;
  wire  T_720;
  wire  T_721;
  wire  T_722;
  wire [7:0] T_723;
  wire [7:0] T_725;
  wire [7:0] T_726;
  wire  T_727;
  wire  T_728;
  wire  T_729;
  wire  T_730;
  wire  T_731;
  wire  T_732;
  wire  T_733;
  wire  T_734;
  wire [7:0] T_738;
  wire [7:0] T_742;
  wire [7:0] T_746;
  wire [7:0] T_750;
  wire [7:0] T_754;
  wire [7:0] T_758;
  wire [7:0] T_762;
  wire [7:0] T_766;
  wire [15:0] T_767;
  wire [15:0] T_768;
  wire [31:0] T_769;
  wire [15:0] T_770;
  wire [15:0] T_771;
  wire [31:0] T_772;
  wire [63:0] T_773;
  wire [63:0] T_774;
  wire [63:0] T_853;
  wire [63:0] T_854;
  wire [63:0] T_855;
  wire  T_859;
  wire [63:0] GEN_2;
  wire [63:0] GEN_7;
  wire [63:0] GEN_8;
  wire  T_865;
  wire  T_867;
  wire  T_868;
  wire [2:0] T_877_0;
  wire [2:0] T_877_1;
  wire [2:0] T_895_0;
  wire [2:0] T_895_1;
  wire [63:0] T_1064;
  wire [63:0] T_1065;
  wire [63:0] GEN_10;
  wire [63:0] GEN_15;
  wire [63:0] GEN_16;
  wire  T_1077;
  wire  T_1078;
  wire [2:0] T_1087_0;
  wire [2:0] T_1087_1;
  wire [2:0] T_1105_0;
  wire [2:0] T_1105_1;
  wire [63:0] GEN_25;
  wire [63:0] T_1274;
  wire [63:0] T_1275;
  wire [63:0] GEN_18;
  wire [63:0] T_1286;
  wire [63:0] GEN_23;
  wire [63:0] GEN_24;
  wire  T_1287;
  wire  T_1288;
  wire  GEN_1;
  reg [31:0] GEN_6;
  Queue_12 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_636_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_636_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_636_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_636_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_636_g_type;
  assign io_tl_grant_bits_data = T_636_data;
  assign io_tiles_0_reset = GEN_1;
  assign io_tiles_0_id = 1'h0;
  assign io_tiles_0_interrupts_meip = io_interrupts_0_meip;
  assign io_tiles_0_interrupts_seip = io_interrupts_0_seip;
  assign io_tiles_0_interrupts_debug = io_interrupts_0_debug;
  assign io_tiles_0_interrupts_mtip = T_1288;
  assign io_tiles_0_interrupts_msip = T_1287;
  assign T_525 = time$ + 64'h1;
  assign T_526 = T_525[63:0];
  assign GEN_0 = io_rtcTick ? T_526 : time$;
  assign T_533_0 = 32'h0;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_568_0 = 3'h0;
  assign T_568_1 = 3'h4;
  assign T_570 = acq_io_deq_bits_a_type == T_568_0;
  assign T_571 = acq_io_deq_bits_a_type == T_568_1;
  assign T_572 = T_570 | T_571;
  assign T_573 = acq_io_deq_bits_is_builtin_type & T_572;
  assign T_574 = acq_io_deq_bits_union[10:8];
  assign T_576 = T_573 ? T_574 : 3'h0;
  assign T_577 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_578 = {T_577,T_576};
  assign addr = T_578[15:0];
  assign rdata = GEN_24;
  assign T_598 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_599 = T_598 ? 3'h1 : 3'h3;
  assign T_600 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_601 = T_600 ? 3'h1 : T_599;
  assign T_602 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_603 = T_602 ? 3'h4 : T_601;
  assign T_604 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_605 = T_604 ? 3'h3 : T_603;
  assign T_606 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_607 = T_606 ? 3'h3 : T_605;
  assign T_608 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_609 = T_608 ? 3'h5 : T_607;
  assign T_610 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_611 = T_610 ? 3'h4 : T_609;
  assign T_636_addr_beat = 3'h0;
  assign T_636_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_636_manager_xact_id = 1'h0;
  assign T_636_is_builtin_type = 1'h1;
  assign T_636_g_type = {{1'd0}, T_611};
  assign T_636_data = rdata;
  assign T_658 = addr[15];
  assign T_659 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_667_0 = 3'h0;
  assign T_667_1 = 3'h4;
  assign T_685_0 = 3'h0;
  assign T_685_1 = 3'h4;
  assign T_697 = acq_io_deq_bits_a_type == 3'h4;
  assign T_698 = acq_io_deq_bits_is_builtin_type & T_697;
  assign T_717 = acq_io_deq_bits_a_type == 3'h3;
  assign T_718 = acq_io_deq_bits_is_builtin_type & T_717;
  assign T_720 = acq_io_deq_bits_a_type == 3'h2;
  assign T_721 = acq_io_deq_bits_is_builtin_type & T_720;
  assign T_722 = T_718 | T_721;
  assign T_723 = acq_io_deq_bits_union[8:1];
  assign T_725 = T_722 ? T_723 : 8'h0;
  assign T_726 = T_698 ? 8'hff : T_725;
  assign T_727 = T_726[0];
  assign T_728 = T_726[1];
  assign T_729 = T_726[2];
  assign T_730 = T_726[3];
  assign T_731 = T_726[4];
  assign T_732 = T_726[5];
  assign T_733 = T_726[6];
  assign T_734 = T_726[7];
  assign T_738 = T_727 ? 8'hff : 8'h0;
  assign T_742 = T_728 ? 8'hff : 8'h0;
  assign T_746 = T_729 ? 8'hff : 8'h0;
  assign T_750 = T_730 ? 8'hff : 8'h0;
  assign T_754 = T_731 ? 8'hff : 8'h0;
  assign T_758 = T_732 ? 8'hff : 8'h0;
  assign T_762 = T_733 ? 8'hff : 8'h0;
  assign T_766 = T_734 ? 8'hff : 8'h0;
  assign T_767 = {T_742,T_738};
  assign T_768 = {T_750,T_746};
  assign T_769 = {T_768,T_767};
  assign T_770 = {T_758,T_754};
  assign T_771 = {T_766,T_762};
  assign T_772 = {T_771,T_770};
  assign T_773 = {T_772,T_769};
  assign T_774 = acq_io_deq_bits_data & T_773;
  assign T_853 = ~ T_773;
  assign T_854 = time$ & T_853;
  assign T_855 = T_774 | T_854;
  assign T_859 = T_659 & T_721;
  assign GEN_2 = T_859 ? T_855 : GEN_0;
  assign GEN_7 = T_658 ? GEN_2 : GEN_0;
  assign GEN_8 = T_658 ? time$ : 64'h0;
  assign T_865 = addr >= 16'h4000;
  assign T_867 = T_658 == 1'h0;
  assign T_868 = T_867 & T_865;
  assign T_877_0 = 3'h0;
  assign T_877_1 = 3'h4;
  assign T_895_0 = 3'h0;
  assign T_895_1 = 3'h4;
  assign T_1064 = timecmp_0 & T_853;
  assign T_1065 = T_774 | T_1064;
  assign GEN_10 = T_859 ? T_1065 : timecmp_0;
  assign GEN_15 = T_868 ? GEN_10 : timecmp_0;
  assign GEN_16 = T_868 ? timecmp_0 : GEN_8;
  assign T_1077 = T_865 == 1'h0;
  assign T_1078 = T_867 & T_1077;
  assign T_1087_0 = 3'h0;
  assign T_1087_1 = 3'h4;
  assign T_1105_0 = 3'h0;
  assign T_1105_1 = 3'h4;
  assign GEN_25 = {{32'd0}, ipi_0};
  assign T_1274 = GEN_25 & T_853;
  assign T_1275 = T_774 | T_1274;
  assign GEN_18 = T_859 ? T_1275 : {{32'd0}, ipi_0};
  assign T_1286 = GEN_25 & 64'h100000001;
  assign GEN_23 = T_1078 ? GEN_18 : {{32'd0}, ipi_0};
  assign GEN_24 = T_1078 ? T_1286 : GEN_16;
  assign T_1287 = ipi_0[0];
  assign T_1288 = time$ >= timecmp_0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_6[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {2{$random}};
  timecmp_0 = GEN_3[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {2{$random}};
  time$ = GEN_4[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  ipi_0 = GEN_5[31:0];
  `endif
  GEN_6 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_868) begin
        if(T_859) begin
          timecmp_0 <= T_1065;
        end
      end
    end
    if(reset) begin
      time$ <= 64'h0;
    end else begin
      if(T_658) begin
        if(T_859) begin
          time$ <= T_855;
        end else begin
          if(io_rtcTick) begin
            time$ <= T_526;
          end
        end
      end else begin
        if(io_rtcTick) begin
          time$ <= T_526;
        end
      end
    end
    if(reset) begin
      ipi_0 <= T_533_0;
    end else begin
      ipi_0 <= GEN_23[31:0];
    end
  end
endmodule
module ROMSlave(
  input   clk,
  input   reset,
  output  io_acquire_ready,
  input   io_acquire_valid,
  input  [25:0] io_acquire_bits_addr_block,
  input  [1:0] io_acquire_bits_client_xact_id,
  input  [2:0] io_acquire_bits_addr_beat,
  input   io_acquire_bits_is_builtin_type,
  input  [2:0] io_acquire_bits_a_type,
  input  [10:0] io_acquire_bits_union,
  input  [63:0] io_acquire_bits_data,
  input   io_grant_ready,
  output  io_grant_valid,
  output [2:0] io_grant_bits_addr_beat,
  output [1:0] io_grant_bits_client_xact_id,
  output  io_grant_bits_manager_xact_id,
  output  io_grant_bits_is_builtin_type,
  output [3:0] io_grant_bits_g_type,
  output [63:0] io_grant_bits_data
);
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [10:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [10:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_446;
  wire  single_beat;
  wire  T_448;
  wire  multi_beat;
  wire  T_450;
  wire  T_451;
  wire  T_452;
  wire  T_453;
  wire  T_455;
  reg [2:0] addr_beat;
  reg [31:0] GEN_54;
  wire  T_457;
  wire [3:0] T_459;
  wire [2:0] T_460;
  wire [2:0] GEN_1;
  wire  T_461;
  wire [2:0] GEN_2;
  wire [63:0] rom_0;
  wire [63:0] rom_1;
  wire [63:0] rom_2;
  wire [63:0] rom_3;
  wire [63:0] rom_4;
  wire [63:0] rom_5;
  wire [63:0] rom_6;
  wire [63:0] rom_7;
  wire [63:0] rom_8;
  wire [63:0] rom_9;
  wire [63:0] rom_10;
  wire [63:0] rom_11;
  wire [63:0] rom_12;
  wire [63:0] rom_13;
  wire [63:0] rom_14;
  wire [63:0] rom_15;
  wire [63:0] rom_16;
  wire [63:0] rom_17;
  wire [63:0] rom_18;
  wire [63:0] rom_19;
  wire [63:0] rom_20;
  wire [63:0] rom_21;
  wire [63:0] rom_22;
  wire [63:0] rom_23;
  wire [63:0] rom_24;
  wire [63:0] rom_25;
  wire [63:0] rom_26;
  wire [63:0] rom_27;
  wire [63:0] rom_28;
  wire [63:0] rom_29;
  wire [63:0] rom_30;
  wire [63:0] rom_31;
  wire [63:0] rom_32;
  wire [63:0] rom_33;
  wire [63:0] rom_34;
  wire [63:0] rom_35;
  wire [63:0] rom_36;
  wire [63:0] rom_37;
  wire [63:0] rom_38;
  wire [63:0] rom_39;
  wire [63:0] rom_40;
  wire [63:0] rom_41;
  wire [63:0] rom_42;
  wire [63:0] rom_43;
  wire [63:0] rom_44;
  wire [63:0] rom_45;
  wire [63:0] rom_46;
  wire [63:0] rom_47;
  wire [63:0] rom_48;
  wire [63:0] rom_49;
  wire [63:0] rom_50;
  wire [63:0] rom_51;
  wire [28:0] raddr;
  wire [5:0] T_520;
  wire  T_522;
  wire  T_524;
  wire  last;
  wire  T_525;
  wire  T_542;
  wire [2:0] T_543;
  wire  T_544;
  wire [2:0] T_545;
  wire  T_546;
  wire [2:0] T_547;
  wire  T_548;
  wire [2:0] T_549;
  wire  T_550;
  wire [2:0] T_551;
  wire  T_552;
  wire [2:0] T_553;
  wire  T_554;
  wire [2:0] T_555;
  wire [2:0] T_579_addr_beat;
  wire [1:0] T_579_client_xact_id;
  wire  T_579_manager_xact_id;
  wire  T_579_is_builtin_type;
  wire [3:0] T_579_g_type;
  wire [63:0] T_579_data;
  wire [63:0] GEN_0;
  wire [63:0] GEN_3;
  wire [63:0] GEN_4;
  wire [63:0] GEN_5;
  wire [63:0] GEN_6;
  wire [63:0] GEN_7;
  wire [63:0] GEN_8;
  wire [63:0] GEN_9;
  wire [63:0] GEN_10;
  wire [63:0] GEN_11;
  wire [63:0] GEN_12;
  wire [63:0] GEN_13;
  wire [63:0] GEN_14;
  wire [63:0] GEN_15;
  wire [63:0] GEN_16;
  wire [63:0] GEN_17;
  wire [63:0] GEN_18;
  wire [63:0] GEN_19;
  wire [63:0] GEN_20;
  wire [63:0] GEN_21;
  wire [63:0] GEN_22;
  wire [63:0] GEN_23;
  wire [63:0] GEN_24;
  wire [63:0] GEN_25;
  wire [63:0] GEN_26;
  wire [63:0] GEN_27;
  wire [63:0] GEN_28;
  wire [63:0] GEN_29;
  wire [63:0] GEN_30;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  wire [63:0] GEN_36;
  wire [63:0] GEN_37;
  wire [63:0] GEN_38;
  wire [63:0] GEN_39;
  wire [63:0] GEN_40;
  wire [63:0] GEN_41;
  wire [63:0] GEN_42;
  wire [63:0] GEN_43;
  wire [63:0] GEN_44;
  wire [63:0] GEN_45;
  wire [63:0] GEN_46;
  wire [63:0] GEN_47;
  wire [63:0] GEN_48;
  wire [63:0] GEN_49;
  wire [63:0] GEN_50;
  wire [63:0] GEN_51;
  wire [63:0] GEN_52;
  wire [63:0] GEN_53;
  Queue_12 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_acquire_ready = acq_io_enq_ready;
  assign io_grant_valid = acq_io_deq_valid;
  assign io_grant_bits_addr_beat = T_579_addr_beat;
  assign io_grant_bits_client_xact_id = T_579_client_xact_id;
  assign io_grant_bits_manager_xact_id = T_579_manager_xact_id;
  assign io_grant_bits_is_builtin_type = T_579_is_builtin_type;
  assign io_grant_bits_g_type = T_579_g_type;
  assign io_grant_bits_data = T_579_data;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_acquire_bits_union;
  assign acq_io_enq_bits_data = io_acquire_bits_data;
  assign acq_io_deq_ready = T_525;
  assign T_446 = acq_io_deq_bits_a_type == 3'h0;
  assign single_beat = acq_io_deq_bits_is_builtin_type & T_446;
  assign T_448 = acq_io_deq_bits_a_type == 3'h1;
  assign multi_beat = acq_io_deq_bits_is_builtin_type & T_448;
  assign T_450 = acq_io_deq_valid == 1'h0;
  assign T_451 = T_450 | single_beat;
  assign T_452 = T_451 | multi_beat;
  assign T_453 = T_452 | reset;
  assign T_455 = T_453 == 1'h0;
  assign T_457 = io_grant_ready & io_grant_valid;
  assign T_459 = addr_beat + 3'h1;
  assign T_460 = T_459[2:0];
  assign GEN_1 = T_457 ? T_460 : addr_beat;
  assign T_461 = io_acquire_ready & io_acquire_valid;
  assign GEN_2 = T_461 ? io_acquire_bits_addr_beat : GEN_1;
  assign rom_0 = 64'h6f;
  assign rom_1 = 64'h102000000000;
  assign rom_2 = 64'h0;
  assign rom_3 = 64'h0;
  assign rom_4 = 64'h200a7b2063696c70;
  assign rom_5 = 64'h7469726f69727020;
  assign rom_6 = 64'h3030303478302079;
  assign rom_7 = 64'h20200a3b30303030;
  assign rom_8 = 64'h20676e69646e6570;
  assign rom_9 = 64'h3031303030347830;
  assign rom_10 = 64'h646e20200a3b3030;
  assign rom_11 = 64'h7d0a3b3220737665;
  assign rom_12 = 64'ha7b206374720a3b;
  assign rom_13 = 64'h3020726464612020;
  assign rom_14 = 64'h6666623030343478;
  assign rom_15 = 64'h61720a3b7d0a3b38;
  assign rom_16 = 64'h203020200a7b206d;
  assign rom_17 = 64'h6461202020200a7b;
  assign rom_18 = 64'h3030387830207264;
  assign rom_19 = 64'h200a3b3030303030;
  assign rom_20 = 64'h20657a6973202020;
  assign rom_21 = 64'h3030303030317830;
  assign rom_22 = 64'h3b7d20200a3b3030;
  assign rom_23 = 64'h65726f630a3b7d0a;
  assign rom_24 = 64'h7b203020200a7b20;
  assign rom_25 = 64'h7b2030202020200a;
  assign rom_26 = 64'h692020202020200a;
  assign rom_27 = 64'h6934367672206173;
  assign rom_28 = 64'h202020200a3b616d;
  assign rom_29 = 64'h6d63656d69742020;
  assign rom_30 = 64'h3030343478302070;
  assign rom_31 = 64'h20200a3b30303034;
  assign rom_32 = 64'h2069706920202020;
  assign rom_33 = 64'h3030303034347830;
  assign rom_34 = 64'h202020200a3b3030;
  assign rom_35 = 64'h7b2063696c702020;
  assign rom_36 = 64'h202020202020200a;
  assign rom_37 = 64'h2020200a7b206d20;
  assign rom_38 = 64'h6569202020202020;
  assign rom_39 = 64'h3230303034783020;
  assign rom_40 = 64'h2020200a3b303030;
  assign rom_41 = 64'h6874202020202020;
  assign rom_42 = 64'h3478302068736572;
  assign rom_43 = 64'h3b30303030303230;
  assign rom_44 = 64'h202020202020200a;
  assign rom_45 = 64'h206d69616c632020;
  assign rom_46 = 64'h3030303230347830;
  assign rom_47 = 64'h202020200a3b3430;
  assign rom_48 = 64'h200a3b7d20202020;
  assign rom_49 = 64'ha3b7d2020202020;
  assign rom_50 = 64'h200a3b7d20202020;
  assign rom_51 = 64'ha3b7d0a3b7d20;
  assign raddr = {acq_io_deq_bits_addr_block,addr_beat};
  assign T_520 = raddr[5:0];
  assign T_522 = multi_beat == 1'h0;
  assign T_524 = addr_beat == 3'h7;
  assign last = T_522 | T_524;
  assign T_525 = io_grant_ready & last;
  assign T_542 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_543 = T_542 ? 3'h1 : 3'h3;
  assign T_544 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_545 = T_544 ? 3'h1 : T_543;
  assign T_546 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_547 = T_546 ? 3'h4 : T_545;
  assign T_548 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_549 = T_548 ? 3'h3 : T_547;
  assign T_550 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_551 = T_550 ? 3'h3 : T_549;
  assign T_552 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_553 = T_552 ? 3'h5 : T_551;
  assign T_554 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_555 = T_554 ? 3'h4 : T_553;
  assign T_579_addr_beat = addr_beat;
  assign T_579_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_579_manager_xact_id = 1'h0;
  assign T_579_is_builtin_type = 1'h1;
  assign T_579_g_type = {{1'd0}, T_555};
  assign T_579_data = GEN_0;
  assign GEN_0 = GEN_53;
  assign GEN_3 = 6'h1 == T_520 ? rom_1 : rom_0;
  assign GEN_4 = 6'h2 == T_520 ? rom_2 : GEN_3;
  assign GEN_5 = 6'h3 == T_520 ? rom_3 : GEN_4;
  assign GEN_6 = 6'h4 == T_520 ? rom_4 : GEN_5;
  assign GEN_7 = 6'h5 == T_520 ? rom_5 : GEN_6;
  assign GEN_8 = 6'h6 == T_520 ? rom_6 : GEN_7;
  assign GEN_9 = 6'h7 == T_520 ? rom_7 : GEN_8;
  assign GEN_10 = 6'h8 == T_520 ? rom_8 : GEN_9;
  assign GEN_11 = 6'h9 == T_520 ? rom_9 : GEN_10;
  assign GEN_12 = 6'ha == T_520 ? rom_10 : GEN_11;
  assign GEN_13 = 6'hb == T_520 ? rom_11 : GEN_12;
  assign GEN_14 = 6'hc == T_520 ? rom_12 : GEN_13;
  assign GEN_15 = 6'hd == T_520 ? rom_13 : GEN_14;
  assign GEN_16 = 6'he == T_520 ? rom_14 : GEN_15;
  assign GEN_17 = 6'hf == T_520 ? rom_15 : GEN_16;
  assign GEN_18 = 6'h10 == T_520 ? rom_16 : GEN_17;
  assign GEN_19 = 6'h11 == T_520 ? rom_17 : GEN_18;
  assign GEN_20 = 6'h12 == T_520 ? rom_18 : GEN_19;
  assign GEN_21 = 6'h13 == T_520 ? rom_19 : GEN_20;
  assign GEN_22 = 6'h14 == T_520 ? rom_20 : GEN_21;
  assign GEN_23 = 6'h15 == T_520 ? rom_21 : GEN_22;
  assign GEN_24 = 6'h16 == T_520 ? rom_22 : GEN_23;
  assign GEN_25 = 6'h17 == T_520 ? rom_23 : GEN_24;
  assign GEN_26 = 6'h18 == T_520 ? rom_24 : GEN_25;
  assign GEN_27 = 6'h19 == T_520 ? rom_25 : GEN_26;
  assign GEN_28 = 6'h1a == T_520 ? rom_26 : GEN_27;
  assign GEN_29 = 6'h1b == T_520 ? rom_27 : GEN_28;
  assign GEN_30 = 6'h1c == T_520 ? rom_28 : GEN_29;
  assign GEN_31 = 6'h1d == T_520 ? rom_29 : GEN_30;
  assign GEN_32 = 6'h1e == T_520 ? rom_30 : GEN_31;
  assign GEN_33 = 6'h1f == T_520 ? rom_31 : GEN_32;
  assign GEN_34 = 6'h20 == T_520 ? rom_32 : GEN_33;
  assign GEN_35 = 6'h21 == T_520 ? rom_33 : GEN_34;
  assign GEN_36 = 6'h22 == T_520 ? rom_34 : GEN_35;
  assign GEN_37 = 6'h23 == T_520 ? rom_35 : GEN_36;
  assign GEN_38 = 6'h24 == T_520 ? rom_36 : GEN_37;
  assign GEN_39 = 6'h25 == T_520 ? rom_37 : GEN_38;
  assign GEN_40 = 6'h26 == T_520 ? rom_38 : GEN_39;
  assign GEN_41 = 6'h27 == T_520 ? rom_39 : GEN_40;
  assign GEN_42 = 6'h28 == T_520 ? rom_40 : GEN_41;
  assign GEN_43 = 6'h29 == T_520 ? rom_41 : GEN_42;
  assign GEN_44 = 6'h2a == T_520 ? rom_42 : GEN_43;
  assign GEN_45 = 6'h2b == T_520 ? rom_43 : GEN_44;
  assign GEN_46 = 6'h2c == T_520 ? rom_44 : GEN_45;
  assign GEN_47 = 6'h2d == T_520 ? rom_45 : GEN_46;
  assign GEN_48 = 6'h2e == T_520 ? rom_46 : GEN_47;
  assign GEN_49 = 6'h2f == T_520 ? rom_47 : GEN_48;
  assign GEN_50 = 6'h30 == T_520 ? rom_48 : GEN_49;
  assign GEN_51 = 6'h31 == T_520 ? rom_49 : GEN_50;
  assign GEN_52 = 6'h32 == T_520 ? rom_50 : GEN_51;
  assign GEN_53 = 6'h33 == T_520 ? rom_51 : GEN_52;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {1{$random}};
  addr_beat = GEN_54[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_461) begin
        addr_beat <= io_acquire_bits_addr_beat;
      end else begin
        if(T_457) begin
          addr_beat <= T_460;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_455) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported ROMSlave operation\n    at Rom.scala:17 assert(!acq.valid || single_beat || multi_beat, \"unsupported ROMSlave operation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_455) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module DefaultCoreplex(
  input   clk,
  input   reset,
  input   io_mem_0_acquire_ready,
  output  io_mem_0_acquire_valid,
  output [25:0] io_mem_0_acquire_bits_addr_block,
  output [1:0] io_mem_0_acquire_bits_client_xact_id,
  output [2:0] io_mem_0_acquire_bits_addr_beat,
  output  io_mem_0_acquire_bits_is_builtin_type,
  output [2:0] io_mem_0_acquire_bits_a_type,
  output [10:0] io_mem_0_acquire_bits_union,
  output [63:0] io_mem_0_acquire_bits_data,
  output  io_mem_0_grant_ready,
  input   io_mem_0_grant_valid,
  input  [2:0] io_mem_0_grant_bits_addr_beat,
  input  [1:0] io_mem_0_grant_bits_client_xact_id,
  input   io_mem_0_grant_bits_manager_xact_id,
  input   io_mem_0_grant_bits_is_builtin_type,
  input  [3:0] io_mem_0_grant_bits_g_type,
  input  [63:0] io_mem_0_grant_bits_data,
  input   io_interrupts_0,
  input   io_interrupts_1,
  output  io_debug_req_ready,
  input   io_debug_req_valid,
  input  [4:0] io_debug_req_bits_addr,
  input  [33:0] io_debug_req_bits_data,
  input  [1:0] io_debug_req_bits_op,
  input   io_debug_resp_ready,
  output  io_debug_resp_valid,
  output [33:0] io_debug_resp_bits_data,
  output [1:0] io_debug_resp_bits_resp,
  input   io_rtcTick
);
  wire  tileResets_0;
  wire  tileList_0_clk;
  wire  tileList_0_reset;
  wire  tileList_0_io_cached_0_acquire_ready;
  wire  tileList_0_io_cached_0_acquire_valid;
  wire [25:0] tileList_0_io_cached_0_acquire_bits_addr_block;
  wire  tileList_0_io_cached_0_acquire_bits_client_xact_id;
  wire [2:0] tileList_0_io_cached_0_acquire_bits_addr_beat;
  wire  tileList_0_io_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] tileList_0_io_cached_0_acquire_bits_a_type;
  wire [10:0] tileList_0_io_cached_0_acquire_bits_union;
  wire [63:0] tileList_0_io_cached_0_acquire_bits_data;
  wire  tileList_0_io_cached_0_probe_ready;
  wire  tileList_0_io_cached_0_probe_valid;
  wire [25:0] tileList_0_io_cached_0_probe_bits_addr_block;
  wire [1:0] tileList_0_io_cached_0_probe_bits_p_type;
  wire  tileList_0_io_cached_0_release_ready;
  wire  tileList_0_io_cached_0_release_valid;
  wire [2:0] tileList_0_io_cached_0_release_bits_addr_beat;
  wire [25:0] tileList_0_io_cached_0_release_bits_addr_block;
  wire  tileList_0_io_cached_0_release_bits_client_xact_id;
  wire  tileList_0_io_cached_0_release_bits_voluntary;
  wire [2:0] tileList_0_io_cached_0_release_bits_r_type;
  wire [63:0] tileList_0_io_cached_0_release_bits_data;
  wire  tileList_0_io_cached_0_grant_ready;
  wire  tileList_0_io_cached_0_grant_valid;
  wire [2:0] tileList_0_io_cached_0_grant_bits_addr_beat;
  wire  tileList_0_io_cached_0_grant_bits_client_xact_id;
  wire [1:0] tileList_0_io_cached_0_grant_bits_manager_xact_id;
  wire  tileList_0_io_cached_0_grant_bits_is_builtin_type;
  wire [3:0] tileList_0_io_cached_0_grant_bits_g_type;
  wire [63:0] tileList_0_io_cached_0_grant_bits_data;
  wire  tileList_0_io_cached_0_grant_bits_manager_id;
  wire  tileList_0_io_cached_0_finish_ready;
  wire  tileList_0_io_cached_0_finish_valid;
  wire [1:0] tileList_0_io_cached_0_finish_bits_manager_xact_id;
  wire  tileList_0_io_cached_0_finish_bits_manager_id;
  wire  tileList_0_io_uncached_0_acquire_ready;
  wire  tileList_0_io_uncached_0_acquire_valid;
  wire [25:0] tileList_0_io_uncached_0_acquire_bits_addr_block;
  wire  tileList_0_io_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] tileList_0_io_uncached_0_acquire_bits_addr_beat;
  wire  tileList_0_io_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] tileList_0_io_uncached_0_acquire_bits_a_type;
  wire [10:0] tileList_0_io_uncached_0_acquire_bits_union;
  wire [63:0] tileList_0_io_uncached_0_acquire_bits_data;
  wire  tileList_0_io_uncached_0_grant_ready;
  wire  tileList_0_io_uncached_0_grant_valid;
  wire [2:0] tileList_0_io_uncached_0_grant_bits_addr_beat;
  wire  tileList_0_io_uncached_0_grant_bits_client_xact_id;
  wire [1:0] tileList_0_io_uncached_0_grant_bits_manager_xact_id;
  wire  tileList_0_io_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] tileList_0_io_uncached_0_grant_bits_g_type;
  wire [63:0] tileList_0_io_uncached_0_grant_bits_data;
  wire  tileList_0_io_prci_reset;
  wire  tileList_0_io_prci_id;
  wire  tileList_0_io_prci_interrupts_meip;
  wire  tileList_0_io_prci_interrupts_seip;
  wire  tileList_0_io_prci_interrupts_debug;
  wire  tileList_0_io_prci_interrupts_mtip;
  wire  tileList_0_io_prci_interrupts_msip;
  wire  PortedTileLinkCrossbar_1_clk;
  wire  PortedTileLinkCrossbar_1_reset;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_block;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_a_type;
  wire [10:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_union;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_data;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_probe_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_probe_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_p_type;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_release_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_release_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_beat;
  wire [25:0] PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_block;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_client_xact_id;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_voluntary;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_r_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_data;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_grant_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_grant_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_client_xact_id;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_is_builtin_type;
  wire [3:0] PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_g_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_data;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_id;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_finish_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_finish_valid;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_id;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_block;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_a_type;
  wire [10:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_union;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_data;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_client_xact_id;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_g_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_0_acquire_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_acquire_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_block;
  wire  PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_is_builtin_type;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_a_type;
  wire [10:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_union;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_grant_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_grant_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_grant_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_xact_id;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_0_grant_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_grant_bits_is_builtin_type;
  wire [3:0] PortedTileLinkCrossbar_1_io_managers_0_grant_bits_g_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_0_grant_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_finish_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_finish_valid;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_0_finish_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_probe_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_probe_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_0_probe_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_0_probe_bits_p_type;
  wire  PortedTileLinkCrossbar_1_io_managers_0_probe_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_release_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_release_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_beat;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_block;
  wire  PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_release_bits_voluntary;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_release_bits_r_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_0_release_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_acquire_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_acquire_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_block;
  wire  PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_is_builtin_type;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_a_type;
  wire [10:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_union;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_grant_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_grant_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_grant_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_xact_id;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_1_grant_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_grant_bits_is_builtin_type;
  wire [3:0] PortedTileLinkCrossbar_1_io_managers_1_grant_bits_g_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_1_grant_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_finish_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_finish_valid;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_1_finish_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_probe_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_probe_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_1_probe_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_1_probe_bits_p_type;
  wire  PortedTileLinkCrossbar_1_io_managers_1_probe_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_release_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_release_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_beat;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_block;
  wire  PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_release_bits_voluntary;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_release_bits_r_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_1_release_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_id;
  wire  L2BroadcastHub_1_clk;
  wire  L2BroadcastHub_1_reset;
  wire  L2BroadcastHub_1_io_inner_acquire_ready;
  wire  L2BroadcastHub_1_io_inner_acquire_valid;
  wire [25:0] L2BroadcastHub_1_io_inner_acquire_bits_addr_block;
  wire  L2BroadcastHub_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_1_io_inner_acquire_bits_addr_beat;
  wire  L2BroadcastHub_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] L2BroadcastHub_1_io_inner_acquire_bits_a_type;
  wire [10:0] L2BroadcastHub_1_io_inner_acquire_bits_union;
  wire [63:0] L2BroadcastHub_1_io_inner_acquire_bits_data;
  wire  L2BroadcastHub_1_io_inner_acquire_bits_client_id;
  wire  L2BroadcastHub_1_io_inner_grant_ready;
  wire  L2BroadcastHub_1_io_inner_grant_valid;
  wire [2:0] L2BroadcastHub_1_io_inner_grant_bits_addr_beat;
  wire  L2BroadcastHub_1_io_inner_grant_bits_client_xact_id;
  wire [1:0] L2BroadcastHub_1_io_inner_grant_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] L2BroadcastHub_1_io_inner_grant_bits_g_type;
  wire [63:0] L2BroadcastHub_1_io_inner_grant_bits_data;
  wire  L2BroadcastHub_1_io_inner_grant_bits_client_id;
  wire  L2BroadcastHub_1_io_inner_finish_ready;
  wire  L2BroadcastHub_1_io_inner_finish_valid;
  wire [1:0] L2BroadcastHub_1_io_inner_finish_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_inner_probe_ready;
  wire  L2BroadcastHub_1_io_inner_probe_valid;
  wire [25:0] L2BroadcastHub_1_io_inner_probe_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_inner_probe_bits_p_type;
  wire  L2BroadcastHub_1_io_inner_probe_bits_client_id;
  wire  L2BroadcastHub_1_io_inner_release_ready;
  wire  L2BroadcastHub_1_io_inner_release_valid;
  wire [2:0] L2BroadcastHub_1_io_inner_release_bits_addr_beat;
  wire [25:0] L2BroadcastHub_1_io_inner_release_bits_addr_block;
  wire  L2BroadcastHub_1_io_inner_release_bits_client_xact_id;
  wire  L2BroadcastHub_1_io_inner_release_bits_voluntary;
  wire [2:0] L2BroadcastHub_1_io_inner_release_bits_r_type;
  wire [63:0] L2BroadcastHub_1_io_inner_release_bits_data;
  wire  L2BroadcastHub_1_io_inner_release_bits_client_id;
  wire  L2BroadcastHub_1_io_incoherent_0;
  wire  L2BroadcastHub_1_io_outer_acquire_ready;
  wire  L2BroadcastHub_1_io_outer_acquire_valid;
  wire [25:0] L2BroadcastHub_1_io_outer_acquire_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_1_io_outer_acquire_bits_addr_beat;
  wire  L2BroadcastHub_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] L2BroadcastHub_1_io_outer_acquire_bits_a_type;
  wire [10:0] L2BroadcastHub_1_io_outer_acquire_bits_union;
  wire [63:0] L2BroadcastHub_1_io_outer_acquire_bits_data;
  wire  L2BroadcastHub_1_io_outer_probe_ready;
  wire  L2BroadcastHub_1_io_outer_probe_valid;
  wire [25:0] L2BroadcastHub_1_io_outer_probe_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_outer_probe_bits_p_type;
  wire  L2BroadcastHub_1_io_outer_release_ready;
  wire  L2BroadcastHub_1_io_outer_release_valid;
  wire [2:0] L2BroadcastHub_1_io_outer_release_bits_addr_beat;
  wire [25:0] L2BroadcastHub_1_io_outer_release_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_outer_release_bits_client_xact_id;
  wire  L2BroadcastHub_1_io_outer_release_bits_voluntary;
  wire [2:0] L2BroadcastHub_1_io_outer_release_bits_r_type;
  wire [63:0] L2BroadcastHub_1_io_outer_release_bits_data;
  wire  L2BroadcastHub_1_io_outer_grant_ready;
  wire  L2BroadcastHub_1_io_outer_grant_valid;
  wire [2:0] L2BroadcastHub_1_io_outer_grant_bits_addr_beat;
  wire [1:0] L2BroadcastHub_1_io_outer_grant_bits_client_xact_id;
  wire  L2BroadcastHub_1_io_outer_grant_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] L2BroadcastHub_1_io_outer_grant_bits_g_type;
  wire [63:0] L2BroadcastHub_1_io_outer_grant_bits_data;
  wire  L2BroadcastHub_1_io_outer_grant_bits_manager_id;
  wire  L2BroadcastHub_1_io_outer_finish_ready;
  wire  L2BroadcastHub_1_io_outer_finish_valid;
  wire  L2BroadcastHub_1_io_outer_finish_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_outer_finish_bits_manager_id;
  wire  MMIOTileLinkManager_1_clk;
  wire  MMIOTileLinkManager_1_reset;
  wire  MMIOTileLinkManager_1_io_inner_acquire_ready;
  wire  MMIOTileLinkManager_1_io_inner_acquire_valid;
  wire [25:0] MMIOTileLinkManager_1_io_inner_acquire_bits_addr_block;
  wire  MMIOTileLinkManager_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] MMIOTileLinkManager_1_io_inner_acquire_bits_addr_beat;
  wire  MMIOTileLinkManager_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] MMIOTileLinkManager_1_io_inner_acquire_bits_a_type;
  wire [10:0] MMIOTileLinkManager_1_io_inner_acquire_bits_union;
  wire [63:0] MMIOTileLinkManager_1_io_inner_acquire_bits_data;
  wire  MMIOTileLinkManager_1_io_inner_acquire_bits_client_id;
  wire  MMIOTileLinkManager_1_io_inner_grant_ready;
  wire  MMIOTileLinkManager_1_io_inner_grant_valid;
  wire [2:0] MMIOTileLinkManager_1_io_inner_grant_bits_addr_beat;
  wire  MMIOTileLinkManager_1_io_inner_grant_bits_client_xact_id;
  wire [1:0] MMIOTileLinkManager_1_io_inner_grant_bits_manager_xact_id;
  wire  MMIOTileLinkManager_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] MMIOTileLinkManager_1_io_inner_grant_bits_g_type;
  wire [63:0] MMIOTileLinkManager_1_io_inner_grant_bits_data;
  wire  MMIOTileLinkManager_1_io_inner_grant_bits_client_id;
  wire  MMIOTileLinkManager_1_io_inner_finish_ready;
  wire  MMIOTileLinkManager_1_io_inner_finish_valid;
  wire [1:0] MMIOTileLinkManager_1_io_inner_finish_bits_manager_xact_id;
  wire  MMIOTileLinkManager_1_io_inner_probe_ready;
  wire  MMIOTileLinkManager_1_io_inner_probe_valid;
  wire [25:0] MMIOTileLinkManager_1_io_inner_probe_bits_addr_block;
  wire [1:0] MMIOTileLinkManager_1_io_inner_probe_bits_p_type;
  wire  MMIOTileLinkManager_1_io_inner_probe_bits_client_id;
  wire  MMIOTileLinkManager_1_io_inner_release_ready;
  wire  MMIOTileLinkManager_1_io_inner_release_valid;
  wire [2:0] MMIOTileLinkManager_1_io_inner_release_bits_addr_beat;
  wire [25:0] MMIOTileLinkManager_1_io_inner_release_bits_addr_block;
  wire  MMIOTileLinkManager_1_io_inner_release_bits_client_xact_id;
  wire  MMIOTileLinkManager_1_io_inner_release_bits_voluntary;
  wire [2:0] MMIOTileLinkManager_1_io_inner_release_bits_r_type;
  wire [63:0] MMIOTileLinkManager_1_io_inner_release_bits_data;
  wire  MMIOTileLinkManager_1_io_inner_release_bits_client_id;
  wire  MMIOTileLinkManager_1_io_incoherent_0;
  wire  MMIOTileLinkManager_1_io_outer_acquire_ready;
  wire  MMIOTileLinkManager_1_io_outer_acquire_valid;
  wire [25:0] MMIOTileLinkManager_1_io_outer_acquire_bits_addr_block;
  wire [1:0] MMIOTileLinkManager_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] MMIOTileLinkManager_1_io_outer_acquire_bits_addr_beat;
  wire  MMIOTileLinkManager_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] MMIOTileLinkManager_1_io_outer_acquire_bits_a_type;
  wire [10:0] MMIOTileLinkManager_1_io_outer_acquire_bits_union;
  wire [63:0] MMIOTileLinkManager_1_io_outer_acquire_bits_data;
  wire  MMIOTileLinkManager_1_io_outer_grant_ready;
  wire  MMIOTileLinkManager_1_io_outer_grant_valid;
  wire [2:0] MMIOTileLinkManager_1_io_outer_grant_bits_addr_beat;
  wire [1:0] MMIOTileLinkManager_1_io_outer_grant_bits_client_xact_id;
  wire  MMIOTileLinkManager_1_io_outer_grant_bits_manager_xact_id;
  wire  MMIOTileLinkManager_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] MMIOTileLinkManager_1_io_outer_grant_bits_g_type;
  wire [63:0] MMIOTileLinkManager_1_io_outer_grant_bits_data;
  wire  TileLinkMemoryInterconnect_1_clk;
  wire  TileLinkMemoryInterconnect_1_reset;
  wire  TileLinkMemoryInterconnect_1_io_in_0_acquire_ready;
  wire  TileLinkMemoryInterconnect_1_io_in_0_acquire_valid;
  wire [25:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_a_type;
  wire [10:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_data;
  wire  TileLinkMemoryInterconnect_1_io_in_0_grant_ready;
  wire  TileLinkMemoryInterconnect_1_io_in_0_grant_valid;
  wire [2:0] TileLinkMemoryInterconnect_1_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkMemoryInterconnect_1_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkMemoryInterconnect_1_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkMemoryInterconnect_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkMemoryInterconnect_1_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkMemoryInterconnect_1_io_in_0_grant_bits_data;
  wire  TileLinkMemoryInterconnect_1_io_out_0_acquire_ready;
  wire  TileLinkMemoryInterconnect_1_io_out_0_acquire_valid;
  wire [25:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_a_type;
  wire [10:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_data;
  wire  TileLinkMemoryInterconnect_1_io_out_0_grant_ready;
  wire  TileLinkMemoryInterconnect_1_io_out_0_grant_valid;
  wire [2:0] TileLinkMemoryInterconnect_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkMemoryInterconnect_1_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkMemoryInterconnect_1_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkMemoryInterconnect_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkMemoryInterconnect_1_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkMemoryInterconnect_1_io_out_0_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_clk;
  wire  ClientTileLinkIOUnwrapper_1_reset;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type;
  wire [10:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_probe_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_probe_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_valid;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type;
  wire [10:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_clk;
  wire  ClientTileLinkEnqueuer_1_reset;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type;
  wire [10:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_probe_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_valid;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  wire [10:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_probe_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_valid;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id;
  wire  ClientUncachedTileLinkEnqueuer_1_clk;
  wire  ClientUncachedTileLinkEnqueuer_1_reset;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_ready;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_valid;
  wire [25:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_data;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_grant_ready;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_grant_valid;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  wire [1:0] ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_data;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_ready;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_valid;
  wire [25:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_grant_ready;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_grant_valid;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id;
  wire [1:0] ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_clk;
  wire  TileLinkRecursiveInterconnect_2_reset;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data;
  wire  PLIC_1_clk;
  wire  PLIC_1_reset;
  wire  PLIC_1_io_devices_0_valid;
  wire  PLIC_1_io_devices_0_ready;
  wire  PLIC_1_io_devices_0_complete;
  wire  PLIC_1_io_devices_1_valid;
  wire  PLIC_1_io_devices_1_ready;
  wire  PLIC_1_io_devices_1_complete;
  wire  PLIC_1_io_harts_0;
  wire  PLIC_1_io_tl_acquire_ready;
  wire  PLIC_1_io_tl_acquire_valid;
  wire [25:0] PLIC_1_io_tl_acquire_bits_addr_block;
  wire [1:0] PLIC_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PLIC_1_io_tl_acquire_bits_addr_beat;
  wire  PLIC_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PLIC_1_io_tl_acquire_bits_a_type;
  wire [10:0] PLIC_1_io_tl_acquire_bits_union;
  wire [63:0] PLIC_1_io_tl_acquire_bits_data;
  wire  PLIC_1_io_tl_grant_ready;
  wire  PLIC_1_io_tl_grant_valid;
  wire [2:0] PLIC_1_io_tl_grant_bits_addr_beat;
  wire [1:0] PLIC_1_io_tl_grant_bits_client_xact_id;
  wire  PLIC_1_io_tl_grant_bits_manager_xact_id;
  wire  PLIC_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PLIC_1_io_tl_grant_bits_g_type;
  wire [63:0] PLIC_1_io_tl_grant_bits_data;
  wire  LevelGateway_2_clk;
  wire  LevelGateway_2_reset;
  wire  LevelGateway_2_io_interrupt;
  wire  LevelGateway_2_io_plic_valid;
  wire  LevelGateway_2_io_plic_ready;
  wire  LevelGateway_2_io_plic_complete;
  wire  LevelGateway_1_1_clk;
  wire  LevelGateway_1_1_reset;
  wire  LevelGateway_1_1_io_interrupt;
  wire  LevelGateway_1_1_io_plic_valid;
  wire  LevelGateway_1_1_io_plic_ready;
  wire  LevelGateway_1_1_io_plic_complete;
  wire  DebugModule_1_clk;
  wire  DebugModule_1_reset;
  wire  DebugModule_1_io_db_req_ready;
  wire  DebugModule_1_io_db_req_valid;
  wire [4:0] DebugModule_1_io_db_req_bits_addr;
  wire [33:0] DebugModule_1_io_db_req_bits_data;
  wire [1:0] DebugModule_1_io_db_req_bits_op;
  wire  DebugModule_1_io_db_resp_ready;
  wire  DebugModule_1_io_db_resp_valid;
  wire [33:0] DebugModule_1_io_db_resp_bits_data;
  wire [1:0] DebugModule_1_io_db_resp_bits_resp;
  wire  DebugModule_1_io_debugInterrupts_0;
  wire  DebugModule_1_io_tl_acquire_ready;
  wire  DebugModule_1_io_tl_acquire_valid;
  wire [25:0] DebugModule_1_io_tl_acquire_bits_addr_block;
  wire [1:0] DebugModule_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] DebugModule_1_io_tl_acquire_bits_addr_beat;
  wire  DebugModule_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] DebugModule_1_io_tl_acquire_bits_a_type;
  wire [10:0] DebugModule_1_io_tl_acquire_bits_union;
  wire [63:0] DebugModule_1_io_tl_acquire_bits_data;
  wire  DebugModule_1_io_tl_grant_ready;
  wire  DebugModule_1_io_tl_grant_valid;
  wire [2:0] DebugModule_1_io_tl_grant_bits_addr_beat;
  wire [1:0] DebugModule_1_io_tl_grant_bits_client_xact_id;
  wire  DebugModule_1_io_tl_grant_bits_manager_xact_id;
  wire  DebugModule_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] DebugModule_1_io_tl_grant_bits_g_type;
  wire [63:0] DebugModule_1_io_tl_grant_bits_data;
  wire  DebugModule_1_io_ndreset;
  wire  DebugModule_1_io_fullreset;
  wire  PRCI_1_clk;
  wire  PRCI_1_reset;
  wire  PRCI_1_io_interrupts_0_meip;
  wire  PRCI_1_io_interrupts_0_seip;
  wire  PRCI_1_io_interrupts_0_debug;
  wire  PRCI_1_io_tl_acquire_ready;
  wire  PRCI_1_io_tl_acquire_valid;
  wire [25:0] PRCI_1_io_tl_acquire_bits_addr_block;
  wire [1:0] PRCI_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PRCI_1_io_tl_acquire_bits_addr_beat;
  wire  PRCI_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PRCI_1_io_tl_acquire_bits_a_type;
  wire [10:0] PRCI_1_io_tl_acquire_bits_union;
  wire [63:0] PRCI_1_io_tl_acquire_bits_data;
  wire  PRCI_1_io_tl_grant_ready;
  wire  PRCI_1_io_tl_grant_valid;
  wire [2:0] PRCI_1_io_tl_grant_bits_addr_beat;
  wire [1:0] PRCI_1_io_tl_grant_bits_client_xact_id;
  wire  PRCI_1_io_tl_grant_bits_manager_xact_id;
  wire  PRCI_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PRCI_1_io_tl_grant_bits_g_type;
  wire [63:0] PRCI_1_io_tl_grant_bits_data;
  wire  PRCI_1_io_tiles_0_reset;
  wire  PRCI_1_io_tiles_0_id;
  wire  PRCI_1_io_tiles_0_interrupts_meip;
  wire  PRCI_1_io_tiles_0_interrupts_seip;
  wire  PRCI_1_io_tiles_0_interrupts_debug;
  wire  PRCI_1_io_tiles_0_interrupts_mtip;
  wire  PRCI_1_io_tiles_0_interrupts_msip;
  wire  PRCI_1_io_rtcTick;
  wire  ROMSlave_1_clk;
  wire  ROMSlave_1_reset;
  wire  ROMSlave_1_io_acquire_ready;
  wire  ROMSlave_1_io_acquire_valid;
  wire [25:0] ROMSlave_1_io_acquire_bits_addr_block;
  wire [1:0] ROMSlave_1_io_acquire_bits_client_xact_id;
  wire [2:0] ROMSlave_1_io_acquire_bits_addr_beat;
  wire  ROMSlave_1_io_acquire_bits_is_builtin_type;
  wire [2:0] ROMSlave_1_io_acquire_bits_a_type;
  wire [10:0] ROMSlave_1_io_acquire_bits_union;
  wire [63:0] ROMSlave_1_io_acquire_bits_data;
  wire  ROMSlave_1_io_grant_ready;
  wire  ROMSlave_1_io_grant_valid;
  wire [2:0] ROMSlave_1_io_grant_bits_addr_beat;
  wire [1:0] ROMSlave_1_io_grant_bits_client_xact_id;
  wire  ROMSlave_1_io_grant_bits_manager_xact_id;
  wire  ROMSlave_1_io_grant_bits_is_builtin_type;
  wire [3:0] ROMSlave_1_io_grant_bits_g_type;
  wire [63:0] ROMSlave_1_io_grant_bits_data;
  wire  GEN_0;
  reg [31:0] GEN_2;
  wire  GEN_1;
  reg [31:0] GEN_3;
  RocketTile tileList_0 (
    .clk(tileList_0_clk),
    .reset(tileList_0_reset),
    .io_cached_0_acquire_ready(tileList_0_io_cached_0_acquire_ready),
    .io_cached_0_acquire_valid(tileList_0_io_cached_0_acquire_valid),
    .io_cached_0_acquire_bits_addr_block(tileList_0_io_cached_0_acquire_bits_addr_block),
    .io_cached_0_acquire_bits_client_xact_id(tileList_0_io_cached_0_acquire_bits_client_xact_id),
    .io_cached_0_acquire_bits_addr_beat(tileList_0_io_cached_0_acquire_bits_addr_beat),
    .io_cached_0_acquire_bits_is_builtin_type(tileList_0_io_cached_0_acquire_bits_is_builtin_type),
    .io_cached_0_acquire_bits_a_type(tileList_0_io_cached_0_acquire_bits_a_type),
    .io_cached_0_acquire_bits_union(tileList_0_io_cached_0_acquire_bits_union),
    .io_cached_0_acquire_bits_data(tileList_0_io_cached_0_acquire_bits_data),
    .io_cached_0_probe_ready(tileList_0_io_cached_0_probe_ready),
    .io_cached_0_probe_valid(tileList_0_io_cached_0_probe_valid),
    .io_cached_0_probe_bits_addr_block(tileList_0_io_cached_0_probe_bits_addr_block),
    .io_cached_0_probe_bits_p_type(tileList_0_io_cached_0_probe_bits_p_type),
    .io_cached_0_release_ready(tileList_0_io_cached_0_release_ready),
    .io_cached_0_release_valid(tileList_0_io_cached_0_release_valid),
    .io_cached_0_release_bits_addr_beat(tileList_0_io_cached_0_release_bits_addr_beat),
    .io_cached_0_release_bits_addr_block(tileList_0_io_cached_0_release_bits_addr_block),
    .io_cached_0_release_bits_client_xact_id(tileList_0_io_cached_0_release_bits_client_xact_id),
    .io_cached_0_release_bits_voluntary(tileList_0_io_cached_0_release_bits_voluntary),
    .io_cached_0_release_bits_r_type(tileList_0_io_cached_0_release_bits_r_type),
    .io_cached_0_release_bits_data(tileList_0_io_cached_0_release_bits_data),
    .io_cached_0_grant_ready(tileList_0_io_cached_0_grant_ready),
    .io_cached_0_grant_valid(tileList_0_io_cached_0_grant_valid),
    .io_cached_0_grant_bits_addr_beat(tileList_0_io_cached_0_grant_bits_addr_beat),
    .io_cached_0_grant_bits_client_xact_id(tileList_0_io_cached_0_grant_bits_client_xact_id),
    .io_cached_0_grant_bits_manager_xact_id(tileList_0_io_cached_0_grant_bits_manager_xact_id),
    .io_cached_0_grant_bits_is_builtin_type(tileList_0_io_cached_0_grant_bits_is_builtin_type),
    .io_cached_0_grant_bits_g_type(tileList_0_io_cached_0_grant_bits_g_type),
    .io_cached_0_grant_bits_data(tileList_0_io_cached_0_grant_bits_data),
    .io_cached_0_grant_bits_manager_id(tileList_0_io_cached_0_grant_bits_manager_id),
    .io_cached_0_finish_ready(tileList_0_io_cached_0_finish_ready),
    .io_cached_0_finish_valid(tileList_0_io_cached_0_finish_valid),
    .io_cached_0_finish_bits_manager_xact_id(tileList_0_io_cached_0_finish_bits_manager_xact_id),
    .io_cached_0_finish_bits_manager_id(tileList_0_io_cached_0_finish_bits_manager_id),
    .io_uncached_0_acquire_ready(tileList_0_io_uncached_0_acquire_ready),
    .io_uncached_0_acquire_valid(tileList_0_io_uncached_0_acquire_valid),
    .io_uncached_0_acquire_bits_addr_block(tileList_0_io_uncached_0_acquire_bits_addr_block),
    .io_uncached_0_acquire_bits_client_xact_id(tileList_0_io_uncached_0_acquire_bits_client_xact_id),
    .io_uncached_0_acquire_bits_addr_beat(tileList_0_io_uncached_0_acquire_bits_addr_beat),
    .io_uncached_0_acquire_bits_is_builtin_type(tileList_0_io_uncached_0_acquire_bits_is_builtin_type),
    .io_uncached_0_acquire_bits_a_type(tileList_0_io_uncached_0_acquire_bits_a_type),
    .io_uncached_0_acquire_bits_union(tileList_0_io_uncached_0_acquire_bits_union),
    .io_uncached_0_acquire_bits_data(tileList_0_io_uncached_0_acquire_bits_data),
    .io_uncached_0_grant_ready(tileList_0_io_uncached_0_grant_ready),
    .io_uncached_0_grant_valid(tileList_0_io_uncached_0_grant_valid),
    .io_uncached_0_grant_bits_addr_beat(tileList_0_io_uncached_0_grant_bits_addr_beat),
    .io_uncached_0_grant_bits_client_xact_id(tileList_0_io_uncached_0_grant_bits_client_xact_id),
    .io_uncached_0_grant_bits_manager_xact_id(tileList_0_io_uncached_0_grant_bits_manager_xact_id),
    .io_uncached_0_grant_bits_is_builtin_type(tileList_0_io_uncached_0_grant_bits_is_builtin_type),
    .io_uncached_0_grant_bits_g_type(tileList_0_io_uncached_0_grant_bits_g_type),
    .io_uncached_0_grant_bits_data(tileList_0_io_uncached_0_grant_bits_data),
    .io_prci_reset(tileList_0_io_prci_reset),
    .io_prci_id(tileList_0_io_prci_id),
    .io_prci_interrupts_meip(tileList_0_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(tileList_0_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(tileList_0_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(tileList_0_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(tileList_0_io_prci_interrupts_msip)
  );
  PortedTileLinkCrossbar PortedTileLinkCrossbar_1 (
    .clk(PortedTileLinkCrossbar_1_clk),
    .reset(PortedTileLinkCrossbar_1_reset),
    .io_clients_cached_0_acquire_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_ready),
    .io_clients_cached_0_acquire_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_valid),
    .io_clients_cached_0_acquire_bits_addr_block(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_block),
    .io_clients_cached_0_acquire_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_client_xact_id),
    .io_clients_cached_0_acquire_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_beat),
    .io_clients_cached_0_acquire_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_is_builtin_type),
    .io_clients_cached_0_acquire_bits_a_type(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_a_type),
    .io_clients_cached_0_acquire_bits_union(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_union),
    .io_clients_cached_0_acquire_bits_data(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_data),
    .io_clients_cached_0_probe_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_probe_ready),
    .io_clients_cached_0_probe_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_probe_valid),
    .io_clients_cached_0_probe_bits_addr_block(PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_addr_block),
    .io_clients_cached_0_probe_bits_p_type(PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_p_type),
    .io_clients_cached_0_release_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_release_ready),
    .io_clients_cached_0_release_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_release_valid),
    .io_clients_cached_0_release_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_beat),
    .io_clients_cached_0_release_bits_addr_block(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_block),
    .io_clients_cached_0_release_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_client_xact_id),
    .io_clients_cached_0_release_bits_voluntary(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_voluntary),
    .io_clients_cached_0_release_bits_r_type(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_r_type),
    .io_clients_cached_0_release_bits_data(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_data),
    .io_clients_cached_0_grant_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_ready),
    .io_clients_cached_0_grant_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_valid),
    .io_clients_cached_0_grant_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_addr_beat),
    .io_clients_cached_0_grant_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_client_xact_id),
    .io_clients_cached_0_grant_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_xact_id),
    .io_clients_cached_0_grant_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_is_builtin_type),
    .io_clients_cached_0_grant_bits_g_type(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_g_type),
    .io_clients_cached_0_grant_bits_data(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_data),
    .io_clients_cached_0_grant_bits_manager_id(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_id),
    .io_clients_cached_0_finish_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_finish_ready),
    .io_clients_cached_0_finish_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_finish_valid),
    .io_clients_cached_0_finish_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_xact_id),
    .io_clients_cached_0_finish_bits_manager_id(PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_id),
    .io_clients_uncached_0_acquire_ready(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_ready),
    .io_clients_uncached_0_acquire_valid(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_valid),
    .io_clients_uncached_0_acquire_bits_addr_block(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_block),
    .io_clients_uncached_0_acquire_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_client_xact_id),
    .io_clients_uncached_0_acquire_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_beat),
    .io_clients_uncached_0_acquire_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_is_builtin_type),
    .io_clients_uncached_0_acquire_bits_a_type(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_a_type),
    .io_clients_uncached_0_acquire_bits_union(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_union),
    .io_clients_uncached_0_acquire_bits_data(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_data),
    .io_clients_uncached_0_grant_ready(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_ready),
    .io_clients_uncached_0_grant_valid(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_valid),
    .io_clients_uncached_0_grant_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_addr_beat),
    .io_clients_uncached_0_grant_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_client_xact_id),
    .io_clients_uncached_0_grant_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_manager_xact_id),
    .io_clients_uncached_0_grant_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_is_builtin_type),
    .io_clients_uncached_0_grant_bits_g_type(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_g_type),
    .io_clients_uncached_0_grant_bits_data(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_data),
    .io_managers_0_acquire_ready(PortedTileLinkCrossbar_1_io_managers_0_acquire_ready),
    .io_managers_0_acquire_valid(PortedTileLinkCrossbar_1_io_managers_0_acquire_valid),
    .io_managers_0_acquire_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_block),
    .io_managers_0_acquire_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_xact_id),
    .io_managers_0_acquire_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_beat),
    .io_managers_0_acquire_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_is_builtin_type),
    .io_managers_0_acquire_bits_a_type(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_a_type),
    .io_managers_0_acquire_bits_union(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_union),
    .io_managers_0_acquire_bits_data(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_data),
    .io_managers_0_acquire_bits_client_id(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_id),
    .io_managers_0_grant_ready(PortedTileLinkCrossbar_1_io_managers_0_grant_ready),
    .io_managers_0_grant_valid(PortedTileLinkCrossbar_1_io_managers_0_grant_valid),
    .io_managers_0_grant_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_addr_beat),
    .io_managers_0_grant_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_xact_id),
    .io_managers_0_grant_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_manager_xact_id),
    .io_managers_0_grant_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_is_builtin_type),
    .io_managers_0_grant_bits_g_type(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_g_type),
    .io_managers_0_grant_bits_data(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_data),
    .io_managers_0_grant_bits_client_id(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_id),
    .io_managers_0_finish_ready(PortedTileLinkCrossbar_1_io_managers_0_finish_ready),
    .io_managers_0_finish_valid(PortedTileLinkCrossbar_1_io_managers_0_finish_valid),
    .io_managers_0_finish_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_managers_0_finish_bits_manager_xact_id),
    .io_managers_0_probe_ready(PortedTileLinkCrossbar_1_io_managers_0_probe_ready),
    .io_managers_0_probe_valid(PortedTileLinkCrossbar_1_io_managers_0_probe_valid),
    .io_managers_0_probe_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_0_probe_bits_addr_block),
    .io_managers_0_probe_bits_p_type(PortedTileLinkCrossbar_1_io_managers_0_probe_bits_p_type),
    .io_managers_0_probe_bits_client_id(PortedTileLinkCrossbar_1_io_managers_0_probe_bits_client_id),
    .io_managers_0_release_ready(PortedTileLinkCrossbar_1_io_managers_0_release_ready),
    .io_managers_0_release_valid(PortedTileLinkCrossbar_1_io_managers_0_release_valid),
    .io_managers_0_release_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_beat),
    .io_managers_0_release_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_block),
    .io_managers_0_release_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_xact_id),
    .io_managers_0_release_bits_voluntary(PortedTileLinkCrossbar_1_io_managers_0_release_bits_voluntary),
    .io_managers_0_release_bits_r_type(PortedTileLinkCrossbar_1_io_managers_0_release_bits_r_type),
    .io_managers_0_release_bits_data(PortedTileLinkCrossbar_1_io_managers_0_release_bits_data),
    .io_managers_0_release_bits_client_id(PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_id),
    .io_managers_1_acquire_ready(PortedTileLinkCrossbar_1_io_managers_1_acquire_ready),
    .io_managers_1_acquire_valid(PortedTileLinkCrossbar_1_io_managers_1_acquire_valid),
    .io_managers_1_acquire_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_block),
    .io_managers_1_acquire_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_xact_id),
    .io_managers_1_acquire_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_beat),
    .io_managers_1_acquire_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_is_builtin_type),
    .io_managers_1_acquire_bits_a_type(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_a_type),
    .io_managers_1_acquire_bits_union(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_union),
    .io_managers_1_acquire_bits_data(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_data),
    .io_managers_1_acquire_bits_client_id(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_id),
    .io_managers_1_grant_ready(PortedTileLinkCrossbar_1_io_managers_1_grant_ready),
    .io_managers_1_grant_valid(PortedTileLinkCrossbar_1_io_managers_1_grant_valid),
    .io_managers_1_grant_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_addr_beat),
    .io_managers_1_grant_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_xact_id),
    .io_managers_1_grant_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_manager_xact_id),
    .io_managers_1_grant_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_is_builtin_type),
    .io_managers_1_grant_bits_g_type(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_g_type),
    .io_managers_1_grant_bits_data(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_data),
    .io_managers_1_grant_bits_client_id(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_id),
    .io_managers_1_finish_ready(PortedTileLinkCrossbar_1_io_managers_1_finish_ready),
    .io_managers_1_finish_valid(PortedTileLinkCrossbar_1_io_managers_1_finish_valid),
    .io_managers_1_finish_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_managers_1_finish_bits_manager_xact_id),
    .io_managers_1_probe_ready(PortedTileLinkCrossbar_1_io_managers_1_probe_ready),
    .io_managers_1_probe_valid(PortedTileLinkCrossbar_1_io_managers_1_probe_valid),
    .io_managers_1_probe_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_1_probe_bits_addr_block),
    .io_managers_1_probe_bits_p_type(PortedTileLinkCrossbar_1_io_managers_1_probe_bits_p_type),
    .io_managers_1_probe_bits_client_id(PortedTileLinkCrossbar_1_io_managers_1_probe_bits_client_id),
    .io_managers_1_release_ready(PortedTileLinkCrossbar_1_io_managers_1_release_ready),
    .io_managers_1_release_valid(PortedTileLinkCrossbar_1_io_managers_1_release_valid),
    .io_managers_1_release_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_beat),
    .io_managers_1_release_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_block),
    .io_managers_1_release_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_xact_id),
    .io_managers_1_release_bits_voluntary(PortedTileLinkCrossbar_1_io_managers_1_release_bits_voluntary),
    .io_managers_1_release_bits_r_type(PortedTileLinkCrossbar_1_io_managers_1_release_bits_r_type),
    .io_managers_1_release_bits_data(PortedTileLinkCrossbar_1_io_managers_1_release_bits_data),
    .io_managers_1_release_bits_client_id(PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_id)
  );
  L2BroadcastHub L2BroadcastHub_1 (
    .clk(L2BroadcastHub_1_clk),
    .reset(L2BroadcastHub_1_reset),
    .io_inner_acquire_ready(L2BroadcastHub_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(L2BroadcastHub_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(L2BroadcastHub_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(L2BroadcastHub_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(L2BroadcastHub_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(L2BroadcastHub_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(L2BroadcastHub_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(L2BroadcastHub_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(L2BroadcastHub_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(L2BroadcastHub_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(L2BroadcastHub_1_io_inner_grant_ready),
    .io_inner_grant_valid(L2BroadcastHub_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(L2BroadcastHub_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(L2BroadcastHub_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(L2BroadcastHub_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(L2BroadcastHub_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(L2BroadcastHub_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(L2BroadcastHub_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(L2BroadcastHub_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(L2BroadcastHub_1_io_inner_finish_ready),
    .io_inner_finish_valid(L2BroadcastHub_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(L2BroadcastHub_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(L2BroadcastHub_1_io_inner_probe_ready),
    .io_inner_probe_valid(L2BroadcastHub_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(L2BroadcastHub_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(L2BroadcastHub_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(L2BroadcastHub_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(L2BroadcastHub_1_io_inner_release_ready),
    .io_inner_release_valid(L2BroadcastHub_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(L2BroadcastHub_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(L2BroadcastHub_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(L2BroadcastHub_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(L2BroadcastHub_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(L2BroadcastHub_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(L2BroadcastHub_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(L2BroadcastHub_1_io_inner_release_bits_client_id),
    .io_incoherent_0(L2BroadcastHub_1_io_incoherent_0),
    .io_outer_acquire_ready(L2BroadcastHub_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(L2BroadcastHub_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(L2BroadcastHub_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(L2BroadcastHub_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(L2BroadcastHub_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(L2BroadcastHub_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(L2BroadcastHub_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(L2BroadcastHub_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(L2BroadcastHub_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(L2BroadcastHub_1_io_outer_probe_ready),
    .io_outer_probe_valid(L2BroadcastHub_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(L2BroadcastHub_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(L2BroadcastHub_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(L2BroadcastHub_1_io_outer_release_ready),
    .io_outer_release_valid(L2BroadcastHub_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(L2BroadcastHub_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(L2BroadcastHub_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(L2BroadcastHub_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(L2BroadcastHub_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(L2BroadcastHub_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(L2BroadcastHub_1_io_outer_release_bits_data),
    .io_outer_grant_ready(L2BroadcastHub_1_io_outer_grant_ready),
    .io_outer_grant_valid(L2BroadcastHub_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(L2BroadcastHub_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(L2BroadcastHub_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(L2BroadcastHub_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(L2BroadcastHub_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(L2BroadcastHub_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(L2BroadcastHub_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(L2BroadcastHub_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(L2BroadcastHub_1_io_outer_finish_ready),
    .io_outer_finish_valid(L2BroadcastHub_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(L2BroadcastHub_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(L2BroadcastHub_1_io_outer_finish_bits_manager_id)
  );
  MMIOTileLinkManager MMIOTileLinkManager_1 (
    .clk(MMIOTileLinkManager_1_clk),
    .reset(MMIOTileLinkManager_1_reset),
    .io_inner_acquire_ready(MMIOTileLinkManager_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(MMIOTileLinkManager_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(MMIOTileLinkManager_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(MMIOTileLinkManager_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(MMIOTileLinkManager_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(MMIOTileLinkManager_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(MMIOTileLinkManager_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(MMIOTileLinkManager_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(MMIOTileLinkManager_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(MMIOTileLinkManager_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(MMIOTileLinkManager_1_io_inner_grant_ready),
    .io_inner_grant_valid(MMIOTileLinkManager_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(MMIOTileLinkManager_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(MMIOTileLinkManager_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(MMIOTileLinkManager_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(MMIOTileLinkManager_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(MMIOTileLinkManager_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(MMIOTileLinkManager_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(MMIOTileLinkManager_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(MMIOTileLinkManager_1_io_inner_finish_ready),
    .io_inner_finish_valid(MMIOTileLinkManager_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(MMIOTileLinkManager_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(MMIOTileLinkManager_1_io_inner_probe_ready),
    .io_inner_probe_valid(MMIOTileLinkManager_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(MMIOTileLinkManager_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(MMIOTileLinkManager_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(MMIOTileLinkManager_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(MMIOTileLinkManager_1_io_inner_release_ready),
    .io_inner_release_valid(MMIOTileLinkManager_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(MMIOTileLinkManager_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(MMIOTileLinkManager_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(MMIOTileLinkManager_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(MMIOTileLinkManager_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(MMIOTileLinkManager_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(MMIOTileLinkManager_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(MMIOTileLinkManager_1_io_inner_release_bits_client_id),
    .io_incoherent_0(MMIOTileLinkManager_1_io_incoherent_0),
    .io_outer_acquire_ready(MMIOTileLinkManager_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(MMIOTileLinkManager_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(MMIOTileLinkManager_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(MMIOTileLinkManager_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(MMIOTileLinkManager_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(MMIOTileLinkManager_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(MMIOTileLinkManager_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(MMIOTileLinkManager_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(MMIOTileLinkManager_1_io_outer_acquire_bits_data),
    .io_outer_grant_ready(MMIOTileLinkManager_1_io_outer_grant_ready),
    .io_outer_grant_valid(MMIOTileLinkManager_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(MMIOTileLinkManager_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(MMIOTileLinkManager_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(MMIOTileLinkManager_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(MMIOTileLinkManager_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(MMIOTileLinkManager_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(MMIOTileLinkManager_1_io_outer_grant_bits_data)
  );
  TileLinkMemoryInterconnect TileLinkMemoryInterconnect_1 (
    .clk(TileLinkMemoryInterconnect_1_clk),
    .reset(TileLinkMemoryInterconnect_1_reset),
    .io_in_0_acquire_ready(TileLinkMemoryInterconnect_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkMemoryInterconnect_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkMemoryInterconnect_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkMemoryInterconnect_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkMemoryInterconnect_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkMemoryInterconnect_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkMemoryInterconnect_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkMemoryInterconnect_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_data)
  );
  ClientTileLinkIOUnwrapper ClientTileLinkIOUnwrapper_1 (
    .clk(ClientTileLinkIOUnwrapper_1_clk),
    .reset(ClientTileLinkIOUnwrapper_1_reset),
    .io_in_acquire_ready(ClientTileLinkIOUnwrapper_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientTileLinkIOUnwrapper_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data),
    .io_in_probe_ready(ClientTileLinkIOUnwrapper_1_io_in_probe_ready),
    .io_in_probe_valid(ClientTileLinkIOUnwrapper_1_io_in_probe_valid),
    .io_in_probe_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block),
    .io_in_probe_bits_p_type(ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type),
    .io_in_release_ready(ClientTileLinkIOUnwrapper_1_io_in_release_ready),
    .io_in_release_valid(ClientTileLinkIOUnwrapper_1_io_in_release_valid),
    .io_in_release_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat),
    .io_in_release_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block),
    .io_in_release_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id),
    .io_in_release_bits_voluntary(ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary),
    .io_in_release_bits_r_type(ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type),
    .io_in_release_bits_data(ClientTileLinkIOUnwrapper_1_io_in_release_bits_data),
    .io_in_grant_ready(ClientTileLinkIOUnwrapper_1_io_in_grant_ready),
    .io_in_grant_valid(ClientTileLinkIOUnwrapper_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data),
    .io_in_grant_bits_manager_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id),
    .io_in_finish_ready(ClientTileLinkIOUnwrapper_1_io_in_finish_ready),
    .io_in_finish_valid(ClientTileLinkIOUnwrapper_1_io_in_finish_valid),
    .io_in_finish_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id),
    .io_in_finish_bits_manager_id(ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id),
    .io_out_acquire_ready(ClientTileLinkIOUnwrapper_1_io_out_acquire_ready),
    .io_out_acquire_valid(ClientTileLinkIOUnwrapper_1_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientTileLinkIOUnwrapper_1_io_out_grant_ready),
    .io_out_grant_valid(ClientTileLinkIOUnwrapper_1_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data)
  );
  ClientTileLinkEnqueuer ClientTileLinkEnqueuer_1 (
    .clk(ClientTileLinkEnqueuer_1_clk),
    .reset(ClientTileLinkEnqueuer_1_reset),
    .io_inner_acquire_ready(ClientTileLinkEnqueuer_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(ClientTileLinkEnqueuer_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data),
    .io_inner_probe_ready(ClientTileLinkEnqueuer_1_io_inner_probe_ready),
    .io_inner_probe_valid(ClientTileLinkEnqueuer_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type),
    .io_inner_release_ready(ClientTileLinkEnqueuer_1_io_inner_release_ready),
    .io_inner_release_valid(ClientTileLinkEnqueuer_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(ClientTileLinkEnqueuer_1_io_inner_release_bits_data),
    .io_inner_grant_ready(ClientTileLinkEnqueuer_1_io_inner_grant_ready),
    .io_inner_grant_valid(ClientTileLinkEnqueuer_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(ClientTileLinkEnqueuer_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_manager_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id),
    .io_inner_finish_ready(ClientTileLinkEnqueuer_1_io_inner_finish_ready),
    .io_inner_finish_valid(ClientTileLinkEnqueuer_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_finish_bits_manager_id(ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id),
    .io_outer_acquire_ready(ClientTileLinkEnqueuer_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(ClientTileLinkEnqueuer_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(ClientTileLinkEnqueuer_1_io_outer_probe_ready),
    .io_outer_probe_valid(ClientTileLinkEnqueuer_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(ClientTileLinkEnqueuer_1_io_outer_release_ready),
    .io_outer_release_valid(ClientTileLinkEnqueuer_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(ClientTileLinkEnqueuer_1_io_outer_release_bits_data),
    .io_outer_grant_ready(ClientTileLinkEnqueuer_1_io_outer_grant_ready),
    .io_outer_grant_valid(ClientTileLinkEnqueuer_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(ClientTileLinkEnqueuer_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(ClientTileLinkEnqueuer_1_io_outer_finish_ready),
    .io_outer_finish_valid(ClientTileLinkEnqueuer_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id)
  );
  ClientUncachedTileLinkEnqueuer ClientUncachedTileLinkEnqueuer_1 (
    .clk(ClientUncachedTileLinkEnqueuer_1_clk),
    .reset(ClientUncachedTileLinkEnqueuer_1_reset),
    .io_inner_acquire_ready(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_data),
    .io_inner_grant_ready(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_ready),
    .io_inner_grant_valid(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_data),
    .io_outer_acquire_ready(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_data),
    .io_outer_grant_ready(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_ready),
    .io_outer_grant_valid(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_data)
  );
  TileLinkRecursiveInterconnect TileLinkRecursiveInterconnect_2 (
    .clk(TileLinkRecursiveInterconnect_2_clk),
    .reset(TileLinkRecursiveInterconnect_2_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_2_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_2_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_2_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_2_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_2_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_2_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_2_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_2_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_2_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_2_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data)
  );
  PLIC PLIC_1 (
    .clk(PLIC_1_clk),
    .reset(PLIC_1_reset),
    .io_devices_0_valid(PLIC_1_io_devices_0_valid),
    .io_devices_0_ready(PLIC_1_io_devices_0_ready),
    .io_devices_0_complete(PLIC_1_io_devices_0_complete),
    .io_devices_1_valid(PLIC_1_io_devices_1_valid),
    .io_devices_1_ready(PLIC_1_io_devices_1_ready),
    .io_devices_1_complete(PLIC_1_io_devices_1_complete),
    .io_harts_0(PLIC_1_io_harts_0),
    .io_tl_acquire_ready(PLIC_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(PLIC_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PLIC_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PLIC_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PLIC_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PLIC_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PLIC_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PLIC_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PLIC_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PLIC_1_io_tl_grant_ready),
    .io_tl_grant_valid(PLIC_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PLIC_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PLIC_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PLIC_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PLIC_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PLIC_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PLIC_1_io_tl_grant_bits_data)
  );
  LevelGateway LevelGateway_2 (
    .clk(LevelGateway_2_clk),
    .reset(LevelGateway_2_reset),
    .io_interrupt(LevelGateway_2_io_interrupt),
    .io_plic_valid(LevelGateway_2_io_plic_valid),
    .io_plic_ready(LevelGateway_2_io_plic_ready),
    .io_plic_complete(LevelGateway_2_io_plic_complete)
  );
  LevelGateway LevelGateway_1_1 (
    .clk(LevelGateway_1_1_clk),
    .reset(LevelGateway_1_1_reset),
    .io_interrupt(LevelGateway_1_1_io_interrupt),
    .io_plic_valid(LevelGateway_1_1_io_plic_valid),
    .io_plic_ready(LevelGateway_1_1_io_plic_ready),
    .io_plic_complete(LevelGateway_1_1_io_plic_complete)
  );
  DebugModule DebugModule_1 (
    .clk(DebugModule_1_clk),
    .reset(DebugModule_1_reset),
    .io_db_req_ready(DebugModule_1_io_db_req_ready),
    .io_db_req_valid(DebugModule_1_io_db_req_valid),
    .io_db_req_bits_addr(DebugModule_1_io_db_req_bits_addr),
    .io_db_req_bits_data(DebugModule_1_io_db_req_bits_data),
    .io_db_req_bits_op(DebugModule_1_io_db_req_bits_op),
    .io_db_resp_ready(DebugModule_1_io_db_resp_ready),
    .io_db_resp_valid(DebugModule_1_io_db_resp_valid),
    .io_db_resp_bits_data(DebugModule_1_io_db_resp_bits_data),
    .io_db_resp_bits_resp(DebugModule_1_io_db_resp_bits_resp),
    .io_debugInterrupts_0(DebugModule_1_io_debugInterrupts_0),
    .io_tl_acquire_ready(DebugModule_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(DebugModule_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(DebugModule_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(DebugModule_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(DebugModule_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(DebugModule_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(DebugModule_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(DebugModule_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(DebugModule_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(DebugModule_1_io_tl_grant_ready),
    .io_tl_grant_valid(DebugModule_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(DebugModule_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(DebugModule_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(DebugModule_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(DebugModule_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(DebugModule_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(DebugModule_1_io_tl_grant_bits_data),
    .io_ndreset(DebugModule_1_io_ndreset),
    .io_fullreset(DebugModule_1_io_fullreset)
  );
  PRCI PRCI_1 (
    .clk(PRCI_1_clk),
    .reset(PRCI_1_reset),
    .io_interrupts_0_meip(PRCI_1_io_interrupts_0_meip),
    .io_interrupts_0_seip(PRCI_1_io_interrupts_0_seip),
    .io_interrupts_0_debug(PRCI_1_io_interrupts_0_debug),
    .io_tl_acquire_ready(PRCI_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(PRCI_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PRCI_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PRCI_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PRCI_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PRCI_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PRCI_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PRCI_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PRCI_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PRCI_1_io_tl_grant_ready),
    .io_tl_grant_valid(PRCI_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PRCI_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PRCI_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PRCI_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PRCI_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PRCI_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PRCI_1_io_tl_grant_bits_data),
    .io_tiles_0_reset(PRCI_1_io_tiles_0_reset),
    .io_tiles_0_id(PRCI_1_io_tiles_0_id),
    .io_tiles_0_interrupts_meip(PRCI_1_io_tiles_0_interrupts_meip),
    .io_tiles_0_interrupts_seip(PRCI_1_io_tiles_0_interrupts_seip),
    .io_tiles_0_interrupts_debug(PRCI_1_io_tiles_0_interrupts_debug),
    .io_tiles_0_interrupts_mtip(PRCI_1_io_tiles_0_interrupts_mtip),
    .io_tiles_0_interrupts_msip(PRCI_1_io_tiles_0_interrupts_msip),
    .io_rtcTick(PRCI_1_io_rtcTick)
  );
  ROMSlave ROMSlave_1 (
    .clk(ROMSlave_1_clk),
    .reset(ROMSlave_1_reset),
    .io_acquire_ready(ROMSlave_1_io_acquire_ready),
    .io_acquire_valid(ROMSlave_1_io_acquire_valid),
    .io_acquire_bits_addr_block(ROMSlave_1_io_acquire_bits_addr_block),
    .io_acquire_bits_client_xact_id(ROMSlave_1_io_acquire_bits_client_xact_id),
    .io_acquire_bits_addr_beat(ROMSlave_1_io_acquire_bits_addr_beat),
    .io_acquire_bits_is_builtin_type(ROMSlave_1_io_acquire_bits_is_builtin_type),
    .io_acquire_bits_a_type(ROMSlave_1_io_acquire_bits_a_type),
    .io_acquire_bits_union(ROMSlave_1_io_acquire_bits_union),
    .io_acquire_bits_data(ROMSlave_1_io_acquire_bits_data),
    .io_grant_ready(ROMSlave_1_io_grant_ready),
    .io_grant_valid(ROMSlave_1_io_grant_valid),
    .io_grant_bits_addr_beat(ROMSlave_1_io_grant_bits_addr_beat),
    .io_grant_bits_client_xact_id(ROMSlave_1_io_grant_bits_client_xact_id),
    .io_grant_bits_manager_xact_id(ROMSlave_1_io_grant_bits_manager_xact_id),
    .io_grant_bits_is_builtin_type(ROMSlave_1_io_grant_bits_is_builtin_type),
    .io_grant_bits_g_type(ROMSlave_1_io_grant_bits_g_type),
    .io_grant_bits_data(ROMSlave_1_io_grant_bits_data)
  );
  assign io_mem_0_acquire_valid = TileLinkMemoryInterconnect_1_io_out_0_acquire_valid;
  assign io_mem_0_acquire_bits_addr_block = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_block;
  assign io_mem_0_acquire_bits_client_xact_id = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_client_xact_id;
  assign io_mem_0_acquire_bits_addr_beat = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_beat;
  assign io_mem_0_acquire_bits_is_builtin_type = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_mem_0_acquire_bits_a_type = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_a_type;
  assign io_mem_0_acquire_bits_union = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_union;
  assign io_mem_0_acquire_bits_data = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_data;
  assign io_mem_0_grant_ready = TileLinkMemoryInterconnect_1_io_out_0_grant_ready;
  assign io_debug_req_ready = DebugModule_1_io_db_req_ready;
  assign io_debug_resp_valid = DebugModule_1_io_db_resp_valid;
  assign io_debug_resp_bits_data = DebugModule_1_io_db_resp_bits_data;
  assign io_debug_resp_bits_resp = DebugModule_1_io_db_resp_bits_resp;
  assign tileResets_0 = reset;
  assign tileList_0_clk = clk;
  assign tileList_0_reset = tileResets_0;
  assign tileList_0_io_cached_0_acquire_ready = PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_ready;
  assign tileList_0_io_cached_0_probe_valid = PortedTileLinkCrossbar_1_io_clients_cached_0_probe_valid;
  assign tileList_0_io_cached_0_probe_bits_addr_block = PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_addr_block;
  assign tileList_0_io_cached_0_probe_bits_p_type = PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_p_type;
  assign tileList_0_io_cached_0_release_ready = PortedTileLinkCrossbar_1_io_clients_cached_0_release_ready;
  assign tileList_0_io_cached_0_grant_valid = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_valid;
  assign tileList_0_io_cached_0_grant_bits_addr_beat = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_addr_beat;
  assign tileList_0_io_cached_0_grant_bits_client_xact_id = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_client_xact_id;
  assign tileList_0_io_cached_0_grant_bits_manager_xact_id = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_xact_id;
  assign tileList_0_io_cached_0_grant_bits_is_builtin_type = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_is_builtin_type;
  assign tileList_0_io_cached_0_grant_bits_g_type = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_g_type;
  assign tileList_0_io_cached_0_grant_bits_data = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_data;
  assign tileList_0_io_cached_0_grant_bits_manager_id = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_id;
  assign tileList_0_io_cached_0_finish_ready = PortedTileLinkCrossbar_1_io_clients_cached_0_finish_ready;
  assign tileList_0_io_uncached_0_acquire_ready = PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_ready;
  assign tileList_0_io_uncached_0_grant_valid = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_valid;
  assign tileList_0_io_uncached_0_grant_bits_addr_beat = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_addr_beat;
  assign tileList_0_io_uncached_0_grant_bits_client_xact_id = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_client_xact_id;
  assign tileList_0_io_uncached_0_grant_bits_manager_xact_id = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_manager_xact_id;
  assign tileList_0_io_uncached_0_grant_bits_is_builtin_type = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_is_builtin_type;
  assign tileList_0_io_uncached_0_grant_bits_g_type = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_g_type;
  assign tileList_0_io_uncached_0_grant_bits_data = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_data;
  assign tileList_0_io_prci_reset = PRCI_1_io_tiles_0_reset;
  assign tileList_0_io_prci_id = PRCI_1_io_tiles_0_id;
  assign tileList_0_io_prci_interrupts_meip = PRCI_1_io_tiles_0_interrupts_meip;
  assign tileList_0_io_prci_interrupts_seip = PRCI_1_io_tiles_0_interrupts_seip;
  assign tileList_0_io_prci_interrupts_debug = PRCI_1_io_tiles_0_interrupts_debug;
  assign tileList_0_io_prci_interrupts_mtip = PRCI_1_io_tiles_0_interrupts_mtip;
  assign tileList_0_io_prci_interrupts_msip = PRCI_1_io_tiles_0_interrupts_msip;
  assign PortedTileLinkCrossbar_1_clk = clk;
  assign PortedTileLinkCrossbar_1_reset = reset;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_valid = tileList_0_io_cached_0_acquire_valid;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_block = tileList_0_io_cached_0_acquire_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_client_xact_id = tileList_0_io_cached_0_acquire_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_beat = tileList_0_io_cached_0_acquire_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_is_builtin_type = tileList_0_io_cached_0_acquire_bits_is_builtin_type;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_a_type = tileList_0_io_cached_0_acquire_bits_a_type;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_union = tileList_0_io_cached_0_acquire_bits_union;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_data = tileList_0_io_cached_0_acquire_bits_data;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_probe_ready = tileList_0_io_cached_0_probe_ready;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_valid = tileList_0_io_cached_0_release_valid;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_beat = tileList_0_io_cached_0_release_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_block = tileList_0_io_cached_0_release_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_client_xact_id = tileList_0_io_cached_0_release_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_voluntary = tileList_0_io_cached_0_release_bits_voluntary;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_r_type = tileList_0_io_cached_0_release_bits_r_type;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_data = tileList_0_io_cached_0_release_bits_data;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_grant_ready = tileList_0_io_cached_0_grant_ready;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_finish_valid = tileList_0_io_cached_0_finish_valid;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_xact_id = tileList_0_io_cached_0_finish_bits_manager_xact_id;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_id = tileList_0_io_cached_0_finish_bits_manager_id;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_valid = tileList_0_io_uncached_0_acquire_valid;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_block = tileList_0_io_uncached_0_acquire_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_client_xact_id = tileList_0_io_uncached_0_acquire_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_beat = tileList_0_io_uncached_0_acquire_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_is_builtin_type = tileList_0_io_uncached_0_acquire_bits_is_builtin_type;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_a_type = tileList_0_io_uncached_0_acquire_bits_a_type;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_union = tileList_0_io_uncached_0_acquire_bits_union;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_data = tileList_0_io_uncached_0_acquire_bits_data;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_ready = tileList_0_io_uncached_0_grant_ready;
  assign PortedTileLinkCrossbar_1_io_managers_0_acquire_ready = L2BroadcastHub_1_io_inner_acquire_ready;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_valid = L2BroadcastHub_1_io_inner_grant_valid;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_addr_beat = L2BroadcastHub_1_io_inner_grant_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_xact_id = L2BroadcastHub_1_io_inner_grant_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_manager_xact_id = L2BroadcastHub_1_io_inner_grant_bits_manager_xact_id;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_is_builtin_type = L2BroadcastHub_1_io_inner_grant_bits_is_builtin_type;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_g_type = L2BroadcastHub_1_io_inner_grant_bits_g_type;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_data = L2BroadcastHub_1_io_inner_grant_bits_data;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_id = L2BroadcastHub_1_io_inner_grant_bits_client_id;
  assign PortedTileLinkCrossbar_1_io_managers_0_finish_ready = L2BroadcastHub_1_io_inner_finish_ready;
  assign PortedTileLinkCrossbar_1_io_managers_0_probe_valid = L2BroadcastHub_1_io_inner_probe_valid;
  assign PortedTileLinkCrossbar_1_io_managers_0_probe_bits_addr_block = L2BroadcastHub_1_io_inner_probe_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_managers_0_probe_bits_p_type = L2BroadcastHub_1_io_inner_probe_bits_p_type;
  assign PortedTileLinkCrossbar_1_io_managers_0_probe_bits_client_id = L2BroadcastHub_1_io_inner_probe_bits_client_id;
  assign PortedTileLinkCrossbar_1_io_managers_0_release_ready = L2BroadcastHub_1_io_inner_release_ready;
  assign PortedTileLinkCrossbar_1_io_managers_1_acquire_ready = MMIOTileLinkManager_1_io_inner_acquire_ready;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_valid = MMIOTileLinkManager_1_io_inner_grant_valid;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_addr_beat = MMIOTileLinkManager_1_io_inner_grant_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_xact_id = MMIOTileLinkManager_1_io_inner_grant_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_manager_xact_id = MMIOTileLinkManager_1_io_inner_grant_bits_manager_xact_id;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_is_builtin_type = MMIOTileLinkManager_1_io_inner_grant_bits_is_builtin_type;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_g_type = MMIOTileLinkManager_1_io_inner_grant_bits_g_type;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_data = MMIOTileLinkManager_1_io_inner_grant_bits_data;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_id = MMIOTileLinkManager_1_io_inner_grant_bits_client_id;
  assign PortedTileLinkCrossbar_1_io_managers_1_finish_ready = MMIOTileLinkManager_1_io_inner_finish_ready;
  assign PortedTileLinkCrossbar_1_io_managers_1_probe_valid = MMIOTileLinkManager_1_io_inner_probe_valid;
  assign PortedTileLinkCrossbar_1_io_managers_1_probe_bits_addr_block = MMIOTileLinkManager_1_io_inner_probe_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_managers_1_probe_bits_p_type = MMIOTileLinkManager_1_io_inner_probe_bits_p_type;
  assign PortedTileLinkCrossbar_1_io_managers_1_probe_bits_client_id = MMIOTileLinkManager_1_io_inner_probe_bits_client_id;
  assign PortedTileLinkCrossbar_1_io_managers_1_release_ready = MMIOTileLinkManager_1_io_inner_release_ready;
  assign L2BroadcastHub_1_clk = clk;
  assign L2BroadcastHub_1_reset = reset;
  assign L2BroadcastHub_1_io_inner_acquire_valid = PortedTileLinkCrossbar_1_io_managers_0_acquire_valid;
  assign L2BroadcastHub_1_io_inner_acquire_bits_addr_block = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_block;
  assign L2BroadcastHub_1_io_inner_acquire_bits_client_xact_id = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_xact_id;
  assign L2BroadcastHub_1_io_inner_acquire_bits_addr_beat = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_beat;
  assign L2BroadcastHub_1_io_inner_acquire_bits_is_builtin_type = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_is_builtin_type;
  assign L2BroadcastHub_1_io_inner_acquire_bits_a_type = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_a_type;
  assign L2BroadcastHub_1_io_inner_acquire_bits_union = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_union;
  assign L2BroadcastHub_1_io_inner_acquire_bits_data = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_data;
  assign L2BroadcastHub_1_io_inner_acquire_bits_client_id = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_id;
  assign L2BroadcastHub_1_io_inner_grant_ready = PortedTileLinkCrossbar_1_io_managers_0_grant_ready;
  assign L2BroadcastHub_1_io_inner_finish_valid = PortedTileLinkCrossbar_1_io_managers_0_finish_valid;
  assign L2BroadcastHub_1_io_inner_finish_bits_manager_xact_id = PortedTileLinkCrossbar_1_io_managers_0_finish_bits_manager_xact_id;
  assign L2BroadcastHub_1_io_inner_probe_ready = PortedTileLinkCrossbar_1_io_managers_0_probe_ready;
  assign L2BroadcastHub_1_io_inner_release_valid = PortedTileLinkCrossbar_1_io_managers_0_release_valid;
  assign L2BroadcastHub_1_io_inner_release_bits_addr_beat = PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_beat;
  assign L2BroadcastHub_1_io_inner_release_bits_addr_block = PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_block;
  assign L2BroadcastHub_1_io_inner_release_bits_client_xact_id = PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_xact_id;
  assign L2BroadcastHub_1_io_inner_release_bits_voluntary = PortedTileLinkCrossbar_1_io_managers_0_release_bits_voluntary;
  assign L2BroadcastHub_1_io_inner_release_bits_r_type = PortedTileLinkCrossbar_1_io_managers_0_release_bits_r_type;
  assign L2BroadcastHub_1_io_inner_release_bits_data = PortedTileLinkCrossbar_1_io_managers_0_release_bits_data;
  assign L2BroadcastHub_1_io_inner_release_bits_client_id = PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_id;
  assign L2BroadcastHub_1_io_incoherent_0 = 1'h0;
  assign L2BroadcastHub_1_io_outer_acquire_ready = ClientTileLinkEnqueuer_1_io_inner_acquire_ready;
  assign L2BroadcastHub_1_io_outer_probe_valid = ClientTileLinkEnqueuer_1_io_inner_probe_valid;
  assign L2BroadcastHub_1_io_outer_probe_bits_addr_block = ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block;
  assign L2BroadcastHub_1_io_outer_probe_bits_p_type = ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type;
  assign L2BroadcastHub_1_io_outer_release_ready = ClientTileLinkEnqueuer_1_io_inner_release_ready;
  assign L2BroadcastHub_1_io_outer_grant_valid = ClientTileLinkEnqueuer_1_io_inner_grant_valid;
  assign L2BroadcastHub_1_io_outer_grant_bits_addr_beat = ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  assign L2BroadcastHub_1_io_outer_grant_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  assign L2BroadcastHub_1_io_outer_grant_bits_manager_xact_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  assign L2BroadcastHub_1_io_outer_grant_bits_is_builtin_type = ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  assign L2BroadcastHub_1_io_outer_grant_bits_g_type = ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  assign L2BroadcastHub_1_io_outer_grant_bits_data = ClientTileLinkEnqueuer_1_io_inner_grant_bits_data;
  assign L2BroadcastHub_1_io_outer_grant_bits_manager_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id;
  assign L2BroadcastHub_1_io_outer_finish_ready = ClientTileLinkEnqueuer_1_io_inner_finish_ready;
  assign MMIOTileLinkManager_1_clk = clk;
  assign MMIOTileLinkManager_1_reset = reset;
  assign MMIOTileLinkManager_1_io_inner_acquire_valid = PortedTileLinkCrossbar_1_io_managers_1_acquire_valid;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_addr_block = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_block;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_client_xact_id = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_xact_id;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_addr_beat = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_beat;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_is_builtin_type = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_is_builtin_type;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_a_type = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_a_type;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_union = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_union;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_data = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_data;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_client_id = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_id;
  assign MMIOTileLinkManager_1_io_inner_grant_ready = PortedTileLinkCrossbar_1_io_managers_1_grant_ready;
  assign MMIOTileLinkManager_1_io_inner_finish_valid = PortedTileLinkCrossbar_1_io_managers_1_finish_valid;
  assign MMIOTileLinkManager_1_io_inner_finish_bits_manager_xact_id = PortedTileLinkCrossbar_1_io_managers_1_finish_bits_manager_xact_id;
  assign MMIOTileLinkManager_1_io_inner_probe_ready = PortedTileLinkCrossbar_1_io_managers_1_probe_ready;
  assign MMIOTileLinkManager_1_io_inner_release_valid = PortedTileLinkCrossbar_1_io_managers_1_release_valid;
  assign MMIOTileLinkManager_1_io_inner_release_bits_addr_beat = PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_beat;
  assign MMIOTileLinkManager_1_io_inner_release_bits_addr_block = PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_block;
  assign MMIOTileLinkManager_1_io_inner_release_bits_client_xact_id = PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_xact_id;
  assign MMIOTileLinkManager_1_io_inner_release_bits_voluntary = PortedTileLinkCrossbar_1_io_managers_1_release_bits_voluntary;
  assign MMIOTileLinkManager_1_io_inner_release_bits_r_type = PortedTileLinkCrossbar_1_io_managers_1_release_bits_r_type;
  assign MMIOTileLinkManager_1_io_inner_release_bits_data = PortedTileLinkCrossbar_1_io_managers_1_release_bits_data;
  assign MMIOTileLinkManager_1_io_inner_release_bits_client_id = PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_id;
  assign MMIOTileLinkManager_1_io_incoherent_0 = GEN_0;
  assign MMIOTileLinkManager_1_io_outer_acquire_ready = ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_ready;
  assign MMIOTileLinkManager_1_io_outer_grant_valid = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_valid;
  assign MMIOTileLinkManager_1_io_outer_grant_bits_addr_beat = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  assign MMIOTileLinkManager_1_io_outer_grant_bits_client_xact_id = {{1'd0}, ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id};
  assign MMIOTileLinkManager_1_io_outer_grant_bits_manager_xact_id = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id[0];
  assign MMIOTileLinkManager_1_io_outer_grant_bits_is_builtin_type = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  assign MMIOTileLinkManager_1_io_outer_grant_bits_g_type = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  assign MMIOTileLinkManager_1_io_outer_grant_bits_data = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_data;
  assign TileLinkMemoryInterconnect_1_clk = clk;
  assign TileLinkMemoryInterconnect_1_reset = reset;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_valid = ClientTileLinkIOUnwrapper_1_io_out_acquire_valid;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_block = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_client_xact_id = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_beat = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_is_builtin_type = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_a_type = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_union = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_data = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data;
  assign TileLinkMemoryInterconnect_1_io_in_0_grant_ready = ClientTileLinkIOUnwrapper_1_io_out_grant_ready;
  assign TileLinkMemoryInterconnect_1_io_out_0_acquire_ready = io_mem_0_acquire_ready;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_valid = io_mem_0_grant_valid;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_addr_beat = io_mem_0_grant_bits_addr_beat;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_client_xact_id = io_mem_0_grant_bits_client_xact_id;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_manager_xact_id = io_mem_0_grant_bits_manager_xact_id;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_is_builtin_type = io_mem_0_grant_bits_is_builtin_type;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_g_type = io_mem_0_grant_bits_g_type;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_data = io_mem_0_grant_bits_data;
  assign ClientTileLinkIOUnwrapper_1_clk = clk;
  assign ClientTileLinkIOUnwrapper_1_reset = reset;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_valid = ClientTileLinkEnqueuer_1_io_outer_acquire_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  assign ClientTileLinkIOUnwrapper_1_io_in_probe_ready = ClientTileLinkEnqueuer_1_io_outer_probe_ready;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_valid = ClientTileLinkEnqueuer_1_io_outer_release_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat = ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block = ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary = ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type = ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_data = ClientTileLinkEnqueuer_1_io_outer_release_bits_data;
  assign ClientTileLinkIOUnwrapper_1_io_in_grant_ready = ClientTileLinkEnqueuer_1_io_outer_grant_ready;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_valid = ClientTileLinkEnqueuer_1_io_outer_finish_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id = ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id = ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_acquire_ready = TileLinkMemoryInterconnect_1_io_in_0_acquire_ready;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_valid = TileLinkMemoryInterconnect_1_io_in_0_grant_valid;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_g_type;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_data;
  assign ClientTileLinkEnqueuer_1_clk = clk;
  assign ClientTileLinkEnqueuer_1_reset = reset;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_valid = L2BroadcastHub_1_io_outer_acquire_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block = L2BroadcastHub_1_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id = L2BroadcastHub_1_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat = L2BroadcastHub_1_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type = L2BroadcastHub_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type = L2BroadcastHub_1_io_outer_acquire_bits_a_type;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union = L2BroadcastHub_1_io_outer_acquire_bits_union;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data = L2BroadcastHub_1_io_outer_acquire_bits_data;
  assign ClientTileLinkEnqueuer_1_io_inner_probe_ready = L2BroadcastHub_1_io_outer_probe_ready;
  assign ClientTileLinkEnqueuer_1_io_inner_release_valid = L2BroadcastHub_1_io_outer_release_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat = L2BroadcastHub_1_io_outer_release_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block = L2BroadcastHub_1_io_outer_release_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id = L2BroadcastHub_1_io_outer_release_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary = L2BroadcastHub_1_io_outer_release_bits_voluntary;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type = L2BroadcastHub_1_io_outer_release_bits_r_type;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_data = L2BroadcastHub_1_io_outer_release_bits_data;
  assign ClientTileLinkEnqueuer_1_io_inner_grant_ready = L2BroadcastHub_1_io_outer_grant_ready;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_valid = L2BroadcastHub_1_io_outer_finish_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id = L2BroadcastHub_1_io_outer_finish_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id = L2BroadcastHub_1_io_outer_finish_bits_manager_id;
  assign ClientTileLinkEnqueuer_1_io_outer_acquire_ready = ClientTileLinkIOUnwrapper_1_io_in_acquire_ready;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_valid = ClientTileLinkIOUnwrapper_1_io_in_probe_valid;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block = ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type = ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type;
  assign ClientTileLinkEnqueuer_1_io_outer_release_ready = ClientTileLinkIOUnwrapper_1_io_in_release_ready;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_valid = ClientTileLinkIOUnwrapper_1_io_in_grant_valid;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_data = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id;
  assign ClientTileLinkEnqueuer_1_io_outer_finish_ready = ClientTileLinkIOUnwrapper_1_io_in_finish_ready;
  assign ClientUncachedTileLinkEnqueuer_1_clk = clk;
  assign ClientUncachedTileLinkEnqueuer_1_reset = reset;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_valid = MMIOTileLinkManager_1_io_outer_acquire_valid;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block = MMIOTileLinkManager_1_io_outer_acquire_bits_addr_block;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id = MMIOTileLinkManager_1_io_outer_acquire_bits_client_xact_id[0];
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat = MMIOTileLinkManager_1_io_outer_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type = MMIOTileLinkManager_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_a_type = MMIOTileLinkManager_1_io_outer_acquire_bits_a_type;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_union = MMIOTileLinkManager_1_io_outer_acquire_bits_union;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_data = MMIOTileLinkManager_1_io_outer_acquire_bits_data;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_grant_ready = MMIOTileLinkManager_1_io_outer_grant_ready;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_ready = TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_valid = TileLinkRecursiveInterconnect_2_io_in_0_grant_valid;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id[0];
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id = {{1'd0}, TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id};
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_g_type = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_data = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_clk = clk;
  assign TileLinkRecursiveInterconnect_2_reset = reset;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_valid;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id = {{1'd0}, ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id};
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_in_0_grant_ready = ClientUncachedTileLinkEnqueuer_1_io_outer_grant_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready = DebugModule_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_valid = DebugModule_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat = DebugModule_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id = DebugModule_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id = DebugModule_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type = DebugModule_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type = DebugModule_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data = DebugModule_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready = ROMSlave_1_io_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_valid = ROMSlave_1_io_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat = ROMSlave_1_io_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id = ROMSlave_1_io_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id = ROMSlave_1_io_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type = ROMSlave_1_io_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type = ROMSlave_1_io_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data = ROMSlave_1_io_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready = PLIC_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_valid = PLIC_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat = PLIC_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id = PLIC_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id = PLIC_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type = PLIC_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type = PLIC_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data = PLIC_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready = PRCI_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_valid = PRCI_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat = PRCI_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id = PRCI_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id = PRCI_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type = PRCI_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type = PRCI_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data = PRCI_1_io_tl_grant_bits_data;
  assign PLIC_1_clk = clk;
  assign PLIC_1_reset = reset;
  assign PLIC_1_io_devices_0_valid = LevelGateway_2_io_plic_valid;
  assign PLIC_1_io_devices_1_valid = LevelGateway_1_1_io_plic_valid;
  assign PLIC_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid;
  assign PLIC_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block;
  assign PLIC_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id;
  assign PLIC_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat;
  assign PLIC_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type;
  assign PLIC_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type;
  assign PLIC_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union;
  assign PLIC_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data;
  assign PLIC_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_2_grant_ready;
  assign LevelGateway_2_clk = clk;
  assign LevelGateway_2_reset = reset;
  assign LevelGateway_2_io_interrupt = io_interrupts_0;
  assign LevelGateway_2_io_plic_ready = PLIC_1_io_devices_0_ready;
  assign LevelGateway_2_io_plic_complete = PLIC_1_io_devices_0_complete;
  assign LevelGateway_1_1_clk = clk;
  assign LevelGateway_1_1_reset = reset;
  assign LevelGateway_1_1_io_interrupt = io_interrupts_1;
  assign LevelGateway_1_1_io_plic_ready = PLIC_1_io_devices_1_ready;
  assign LevelGateway_1_1_io_plic_complete = PLIC_1_io_devices_1_complete;
  assign DebugModule_1_clk = clk;
  assign DebugModule_1_reset = reset;
  assign DebugModule_1_io_db_req_valid = io_debug_req_valid;
  assign DebugModule_1_io_db_req_bits_addr = io_debug_req_bits_addr;
  assign DebugModule_1_io_db_req_bits_data = io_debug_req_bits_data;
  assign DebugModule_1_io_db_req_bits_op = io_debug_req_bits_op;
  assign DebugModule_1_io_db_resp_ready = io_debug_resp_ready;
  assign DebugModule_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid;
  assign DebugModule_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block;
  assign DebugModule_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id;
  assign DebugModule_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat;
  assign DebugModule_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type;
  assign DebugModule_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type;
  assign DebugModule_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union;
  assign DebugModule_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data;
  assign DebugModule_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_0_grant_ready;
  assign PRCI_1_clk = clk;
  assign PRCI_1_reset = reset;
  assign PRCI_1_io_interrupts_0_meip = PLIC_1_io_harts_0;
  assign PRCI_1_io_interrupts_0_seip = GEN_1;
  assign PRCI_1_io_interrupts_0_debug = DebugModule_1_io_debugInterrupts_0;
  assign PRCI_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid;
  assign PRCI_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block;
  assign PRCI_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id;
  assign PRCI_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat;
  assign PRCI_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type;
  assign PRCI_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type;
  assign PRCI_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union;
  assign PRCI_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data;
  assign PRCI_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_3_grant_ready;
  assign PRCI_1_io_rtcTick = io_rtcTick;
  assign ROMSlave_1_clk = clk;
  assign ROMSlave_1_reset = reset;
  assign ROMSlave_1_io_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid;
  assign ROMSlave_1_io_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block;
  assign ROMSlave_1_io_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id;
  assign ROMSlave_1_io_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat;
  assign ROMSlave_1_io_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type;
  assign ROMSlave_1_io_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type;
  assign ROMSlave_1_io_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union;
  assign ROMSlave_1_io_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data;
  assign ROMSlave_1_io_grant_ready = TileLinkRecursiveInterconnect_2_io_out_1_grant_ready;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_0 = GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_3[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_2 = {1{$random}};
  GEN_3 = {1{$random}};
  end
`endif
endmodule
module ReorderQueue_2(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_data_addr_beat,
  input   io_enq_bits_data_subblock,
  input  [1:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [1:0] io_deq_tag,
  output [2:0] io_deq_data_addr_beat,
  output  io_deq_data_subblock,
  output  io_deq_matches
);
  reg [2:0] T_229_addr_beat [0:3];
  reg [31:0] GEN_14;
  wire [2:0] T_229_addr_beat_T_245_data;
  wire [1:0] T_229_addr_beat_T_245_addr;
  wire  T_229_addr_beat_T_245_en;
  wire [2:0] T_229_addr_beat_T_271_data;
  wire [1:0] T_229_addr_beat_T_271_addr;
  wire  T_229_addr_beat_T_271_mask;
  wire  T_229_addr_beat_T_271_en;
  reg  T_229_subblock [0:3];
  reg [31:0] GEN_15;
  wire  T_229_subblock_T_245_data;
  wire [1:0] T_229_subblock_T_245_addr;
  wire  T_229_subblock_T_245_en;
  wire  T_229_subblock_T_271_data;
  wire [1:0] T_229_subblock_T_271_addr;
  wire  T_229_subblock_T_271_mask;
  wire  T_229_subblock_T_271_en;
  wire  T_239_0;
  wire  T_239_1;
  wire  T_239_2;
  wire  T_239_3;
  reg  T_243_0;
  reg [31:0] GEN_16;
  reg  T_243_1;
  reg [31:0] GEN_17;
  reg  T_243_2;
  reg [31:0] GEN_18;
  reg  T_243_3;
  reg [31:0] GEN_19;
  wire  GEN_0;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_1;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  T_269;
  wire  T_270;
  wire  GEN_2;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_3;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  assign io_enq_ready = GEN_0;
  assign io_deq_data_addr_beat = T_229_addr_beat_T_245_data;
  assign io_deq_data_subblock = T_229_subblock_T_245_data;
  assign io_deq_matches = T_269;
  assign T_229_addr_beat_T_245_addr = io_deq_tag;
  assign T_229_addr_beat_T_245_en = 1'h1;
  assign T_229_addr_beat_T_245_data = T_229_addr_beat[T_229_addr_beat_T_245_addr];
  assign T_229_addr_beat_T_271_data = io_enq_bits_data_addr_beat;
  assign T_229_addr_beat_T_271_addr = io_enq_bits_tag;
  assign T_229_addr_beat_T_271_mask = T_270;
  assign T_229_addr_beat_T_271_en = T_270;
  assign T_229_subblock_T_245_addr = io_deq_tag;
  assign T_229_subblock_T_245_en = 1'h1;
  assign T_229_subblock_T_245_data = T_229_subblock[T_229_subblock_T_245_addr];
  assign T_229_subblock_T_271_data = io_enq_bits_data_subblock;
  assign T_229_subblock_T_271_addr = io_enq_bits_tag;
  assign T_229_subblock_T_271_mask = T_270;
  assign T_229_subblock_T_271_en = T_270;
  assign T_239_0 = 1'h1;
  assign T_239_1 = 1'h1;
  assign T_239_2 = 1'h1;
  assign T_239_3 = 1'h1;
  assign GEN_0 = GEN_6;
  assign GEN_4 = 2'h1 == io_enq_bits_tag ? T_243_1 : T_243_0;
  assign GEN_5 = 2'h2 == io_enq_bits_tag ? T_243_2 : GEN_4;
  assign GEN_6 = 2'h3 == io_enq_bits_tag ? T_243_3 : GEN_5;
  assign GEN_1 = GEN_9;
  assign GEN_7 = 2'h1 == io_deq_tag ? T_243_1 : T_243_0;
  assign GEN_8 = 2'h2 == io_deq_tag ? T_243_2 : GEN_7;
  assign GEN_9 = 2'h3 == io_deq_tag ? T_243_3 : GEN_8;
  assign T_269 = GEN_1 == 1'h0;
  assign T_270 = io_enq_valid & io_enq_ready;
  assign GEN_2 = 1'h0;
  assign GEN_10 = 2'h0 == io_enq_bits_tag ? GEN_2 : T_243_0;
  assign GEN_11 = 2'h1 == io_enq_bits_tag ? GEN_2 : T_243_1;
  assign GEN_12 = 2'h2 == io_enq_bits_tag ? GEN_2 : T_243_2;
  assign GEN_13 = 2'h3 == io_enq_bits_tag ? GEN_2 : T_243_3;
  assign GEN_22 = T_270 ? GEN_10 : T_243_0;
  assign GEN_23 = T_270 ? GEN_11 : T_243_1;
  assign GEN_24 = T_270 ? GEN_12 : T_243_2;
  assign GEN_25 = T_270 ? GEN_13 : T_243_3;
  assign GEN_3 = 1'h1;
  assign GEN_26 = 2'h0 == io_deq_tag ? GEN_3 : GEN_22;
  assign GEN_27 = 2'h1 == io_deq_tag ? GEN_3 : GEN_23;
  assign GEN_28 = 2'h2 == io_deq_tag ? GEN_3 : GEN_24;
  assign GEN_29 = 2'h3 == io_deq_tag ? GEN_3 : GEN_25;
  assign GEN_31 = io_deq_valid ? GEN_26 : GEN_22;
  assign GEN_32 = io_deq_valid ? GEN_27 : GEN_23;
  assign GEN_33 = io_deq_valid ? GEN_28 : GEN_24;
  assign GEN_34 = io_deq_valid ? GEN_29 : GEN_25;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_14 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    T_229_addr_beat[initvar] = GEN_14[2:0];
  `endif
  GEN_15 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    T_229_subblock[initvar] = GEN_15[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_16 = {1{$random}};
  T_243_0 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {1{$random}};
  T_243_1 = GEN_17[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {1{$random}};
  T_243_2 = GEN_18[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_19 = {1{$random}};
  T_243_3 = GEN_19[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(T_229_addr_beat_T_271_en & T_229_addr_beat_T_271_mask) begin
      T_229_addr_beat[T_229_addr_beat_T_271_addr] <= T_229_addr_beat_T_271_data;
    end
    if(T_229_subblock_T_271_en & T_229_subblock_T_271_mask) begin
      T_229_subblock[T_229_subblock_T_271_addr] <= T_229_subblock_T_271_data;
    end
    if(reset) begin
      T_243_0 <= T_239_0;
    end else begin
      if(io_deq_valid) begin
        if(2'h0 == io_deq_tag) begin
          T_243_0 <= GEN_3;
        end else begin
          if(T_270) begin
            if(2'h0 == io_enq_bits_tag) begin
              T_243_0 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_270) begin
          if(2'h0 == io_enq_bits_tag) begin
            T_243_0 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_243_1 <= T_239_1;
    end else begin
      if(io_deq_valid) begin
        if(2'h1 == io_deq_tag) begin
          T_243_1 <= GEN_3;
        end else begin
          if(T_270) begin
            if(2'h1 == io_enq_bits_tag) begin
              T_243_1 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_270) begin
          if(2'h1 == io_enq_bits_tag) begin
            T_243_1 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_243_2 <= T_239_2;
    end else begin
      if(io_deq_valid) begin
        if(2'h2 == io_deq_tag) begin
          T_243_2 <= GEN_3;
        end else begin
          if(T_270) begin
            if(2'h2 == io_enq_bits_tag) begin
              T_243_2 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_270) begin
          if(2'h2 == io_enq_bits_tag) begin
            T_243_2 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_243_3 <= T_239_3;
    end else begin
      if(io_deq_valid) begin
        if(2'h3 == io_deq_tag) begin
          T_243_3 <= GEN_3;
        end else begin
          if(T_270) begin
            if(2'h3 == io_enq_bits_tag) begin
              T_243_3 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_270) begin
          if(2'h3 == io_enq_bits_tag) begin
            T_243_3 <= GEN_2;
          end
        end
      end
    end
  end
endmodule
module IdMapper(
  input   clk,
  input   reset,
  input   io_req_valid,
  output  io_req_ready,
  input  [1:0] io_req_in_id,
  output [4:0] io_req_out_id,
  input   io_resp_valid,
  output  io_resp_matches,
  input  [4:0] io_resp_out_id,
  output [1:0] io_resp_in_id
);
  assign io_req_ready = 1'h1;
  assign io_req_out_id = {{3'd0}, io_req_in_id};
  assign io_resp_matches = 1'h1;
  assign io_resp_in_id = io_resp_out_id[1:0];
endmodule
module LockingArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire  GEN_0_bits_manager_xact_id;
  wire  GEN_0_bits_is_builtin_type;
  wire [3:0] GEN_0_bits_g_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_0_bits_client_id;
  wire  GEN_8;
  wire  GEN_9;
  wire [2:0] GEN_10;
  wire [1:0] GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire [3:0] GEN_14;
  wire [63:0] GEN_15;
  wire  GEN_16;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire  GEN_1_bits_manager_xact_id;
  wire  GEN_1_bits_is_builtin_type;
  wire [3:0] GEN_1_bits_g_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_1_bits_client_id;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire  GEN_2_bits_manager_xact_id;
  wire  GEN_2_bits_is_builtin_type;
  wire [3:0] GEN_2_bits_g_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_2_bits_client_id;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire  GEN_3_bits_manager_xact_id;
  wire  GEN_3_bits_is_builtin_type;
  wire [3:0] GEN_3_bits_g_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_3_bits_client_id;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire  GEN_4_bits_manager_xact_id;
  wire  GEN_4_bits_is_builtin_type;
  wire [3:0] GEN_4_bits_g_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_4_bits_client_id;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire  GEN_5_bits_manager_xact_id;
  wire  GEN_5_bits_is_builtin_type;
  wire [3:0] GEN_5_bits_g_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_5_bits_client_id;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire  GEN_6_bits_manager_xact_id;
  wire  GEN_6_bits_is_builtin_type;
  wire [3:0] GEN_6_bits_g_type;
  wire [63:0] GEN_6_bits_data;
  wire  GEN_6_bits_client_id;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [2:0] GEN_7_bits_addr_beat;
  wire [1:0] GEN_7_bits_client_xact_id;
  wire  GEN_7_bits_manager_xact_id;
  wire  GEN_7_bits_is_builtin_type;
  wire [3:0] GEN_7_bits_g_type;
  wire [63:0] GEN_7_bits_data;
  wire  GEN_7_bits_client_id;
  reg [2:0] T_766;
  reg [31:0] GEN_1;
  reg  T_768;
  reg [31:0] GEN_2;
  wire  T_770;
  wire [2:0] T_778_0;
  wire [3:0] GEN_0;
  wire  T_780;
  wire  T_781;
  wire  T_782;
  wire  T_784;
  wire  T_785;
  wire [3:0] T_789;
  wire [2:0] T_790;
  wire  GEN_80;
  wire [2:0] GEN_81;
  wire  GEN_82;
  wire  T_793;
  wire  T_795;
  wire  T_796;
  wire  T_797;
  wire  T_800;
  wire  T_801;
  wire  GEN_83;
  assign io_in_0_ready = T_797;
  assign io_in_1_ready = T_801;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = GEN_3_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_g_type = GEN_5_bits_g_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_out_bits_client_id = GEN_7_bits_client_id;
  assign io_chosen = GEN_82;
  assign choice = GEN_83;
  assign GEN_0_ready = GEN_8;
  assign GEN_0_valid = GEN_9;
  assign GEN_0_bits_addr_beat = GEN_10;
  assign GEN_0_bits_client_xact_id = GEN_11;
  assign GEN_0_bits_manager_xact_id = GEN_12;
  assign GEN_0_bits_is_builtin_type = GEN_13;
  assign GEN_0_bits_g_type = GEN_14;
  assign GEN_0_bits_data = GEN_15;
  assign GEN_0_bits_client_id = GEN_16;
  assign GEN_8 = io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_9 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_11 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_13 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_14 = io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_15 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_16 = io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_1_ready = GEN_8;
  assign GEN_1_valid = GEN_9;
  assign GEN_1_bits_addr_beat = GEN_10;
  assign GEN_1_bits_client_xact_id = GEN_11;
  assign GEN_1_bits_manager_xact_id = GEN_12;
  assign GEN_1_bits_is_builtin_type = GEN_13;
  assign GEN_1_bits_g_type = GEN_14;
  assign GEN_1_bits_data = GEN_15;
  assign GEN_1_bits_client_id = GEN_16;
  assign GEN_2_ready = GEN_8;
  assign GEN_2_valid = GEN_9;
  assign GEN_2_bits_addr_beat = GEN_10;
  assign GEN_2_bits_client_xact_id = GEN_11;
  assign GEN_2_bits_manager_xact_id = GEN_12;
  assign GEN_2_bits_is_builtin_type = GEN_13;
  assign GEN_2_bits_g_type = GEN_14;
  assign GEN_2_bits_data = GEN_15;
  assign GEN_2_bits_client_id = GEN_16;
  assign GEN_3_ready = GEN_8;
  assign GEN_3_valid = GEN_9;
  assign GEN_3_bits_addr_beat = GEN_10;
  assign GEN_3_bits_client_xact_id = GEN_11;
  assign GEN_3_bits_manager_xact_id = GEN_12;
  assign GEN_3_bits_is_builtin_type = GEN_13;
  assign GEN_3_bits_g_type = GEN_14;
  assign GEN_3_bits_data = GEN_15;
  assign GEN_3_bits_client_id = GEN_16;
  assign GEN_4_ready = GEN_8;
  assign GEN_4_valid = GEN_9;
  assign GEN_4_bits_addr_beat = GEN_10;
  assign GEN_4_bits_client_xact_id = GEN_11;
  assign GEN_4_bits_manager_xact_id = GEN_12;
  assign GEN_4_bits_is_builtin_type = GEN_13;
  assign GEN_4_bits_g_type = GEN_14;
  assign GEN_4_bits_data = GEN_15;
  assign GEN_4_bits_client_id = GEN_16;
  assign GEN_5_ready = GEN_8;
  assign GEN_5_valid = GEN_9;
  assign GEN_5_bits_addr_beat = GEN_10;
  assign GEN_5_bits_client_xact_id = GEN_11;
  assign GEN_5_bits_manager_xact_id = GEN_12;
  assign GEN_5_bits_is_builtin_type = GEN_13;
  assign GEN_5_bits_g_type = GEN_14;
  assign GEN_5_bits_data = GEN_15;
  assign GEN_5_bits_client_id = GEN_16;
  assign GEN_6_ready = GEN_8;
  assign GEN_6_valid = GEN_9;
  assign GEN_6_bits_addr_beat = GEN_10;
  assign GEN_6_bits_client_xact_id = GEN_11;
  assign GEN_6_bits_manager_xact_id = GEN_12;
  assign GEN_6_bits_is_builtin_type = GEN_13;
  assign GEN_6_bits_g_type = GEN_14;
  assign GEN_6_bits_data = GEN_15;
  assign GEN_6_bits_client_id = GEN_16;
  assign GEN_7_ready = GEN_8;
  assign GEN_7_valid = GEN_9;
  assign GEN_7_bits_addr_beat = GEN_10;
  assign GEN_7_bits_client_xact_id = GEN_11;
  assign GEN_7_bits_manager_xact_id = GEN_12;
  assign GEN_7_bits_is_builtin_type = GEN_13;
  assign GEN_7_bits_g_type = GEN_14;
  assign GEN_7_bits_data = GEN_15;
  assign GEN_7_bits_client_id = GEN_16;
  assign T_770 = T_766 != 3'h0;
  assign T_778_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_778_0};
  assign T_780 = io_out_bits_g_type == GEN_0;
  assign T_781 = io_out_bits_g_type == 4'h0;
  assign T_782 = io_out_bits_is_builtin_type ? T_780 : T_781;
  assign T_784 = io_out_ready & io_out_valid;
  assign T_785 = T_784 & T_782;
  assign T_789 = T_766 + 3'h1;
  assign T_790 = T_789[2:0];
  assign GEN_80 = T_785 ? io_chosen : T_768;
  assign GEN_81 = T_785 ? T_790 : T_766;
  assign GEN_82 = T_770 ? T_768 : choice;
  assign T_793 = io_in_0_valid == 1'h0;
  assign T_795 = T_768 == 1'h0;
  assign T_796 = T_770 ? T_795 : 1'h1;
  assign T_797 = T_796 & io_out_ready;
  assign T_800 = T_770 ? T_768 : T_793;
  assign T_801 = T_800 & io_out_ready;
  assign GEN_83 = io_in_0_valid ? 1'h0 : 1'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_766 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_768 = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_766 <= 3'h0;
    end else begin
      if(T_785) begin
        T_766 <= T_790;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_785) begin
        T_768 <= io_chosen;
      end
    end
  end
endmodule
module NastiIOTileLinkIOConverter(
  input   clk,
  input   reset,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [10:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  input   io_nasti_aw_ready,
  output  io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  output [7:0] io_nasti_aw_bits_len,
  output [2:0] io_nasti_aw_bits_size,
  output [1:0] io_nasti_aw_bits_burst,
  output  io_nasti_aw_bits_lock,
  output [3:0] io_nasti_aw_bits_cache,
  output [2:0] io_nasti_aw_bits_prot,
  output [3:0] io_nasti_aw_bits_qos,
  output [3:0] io_nasti_aw_bits_region,
  output [4:0] io_nasti_aw_bits_id,
  output  io_nasti_aw_bits_user,
  input   io_nasti_w_ready,
  output  io_nasti_w_valid,
  output [63:0] io_nasti_w_bits_data,
  output  io_nasti_w_bits_last,
  output [4:0] io_nasti_w_bits_id,
  output [7:0] io_nasti_w_bits_strb,
  output  io_nasti_w_bits_user,
  output  io_nasti_b_ready,
  input   io_nasti_b_valid,
  input  [1:0] io_nasti_b_bits_resp,
  input  [4:0] io_nasti_b_bits_id,
  input   io_nasti_b_bits_user,
  input   io_nasti_ar_ready,
  output  io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output [7:0] io_nasti_ar_bits_len,
  output [2:0] io_nasti_ar_bits_size,
  output [1:0] io_nasti_ar_bits_burst,
  output  io_nasti_ar_bits_lock,
  output [3:0] io_nasti_ar_bits_cache,
  output [2:0] io_nasti_ar_bits_prot,
  output [3:0] io_nasti_ar_bits_qos,
  output [3:0] io_nasti_ar_bits_region,
  output [4:0] io_nasti_ar_bits_id,
  output  io_nasti_ar_bits_user,
  output  io_nasti_r_ready,
  input   io_nasti_r_valid,
  input  [1:0] io_nasti_r_bits_resp,
  input  [63:0] io_nasti_r_bits_data,
  input   io_nasti_r_bits_last,
  input  [4:0] io_nasti_r_bits_id,
  input   io_nasti_r_bits_user
);
  wire [2:0] T_688_0;
  wire [2:0] T_688_1;
  wire [2:0] T_688_2;
  wire  T_690;
  wire  T_691;
  wire  T_692;
  wire  T_693;
  wire  T_694;
  wire  has_data;
  wire [2:0] T_703_0;
  wire [2:0] T_703_1;
  wire [2:0] T_703_2;
  wire  T_705;
  wire  T_706;
  wire  T_707;
  wire  T_708;
  wire  T_709;
  wire  is_subblock;
  wire [2:0] T_718_0;
  wire  T_720;
  wire  is_multibeat;
  wire  T_721;
  wire  T_722;
  reg [2:0] tl_cnt_out;
  reg [31:0] GEN_11;
  wire  T_725;
  wire [3:0] T_727;
  wire [2:0] T_728;
  wire [2:0] GEN_0;
  wire  tl_wrap_out;
  wire  T_730;
  wire  get_valid;
  wire  put_valid;
  wire  roq_clk;
  wire  roq_reset;
  wire  roq_io_enq_ready;
  wire  roq_io_enq_valid;
  wire [2:0] roq_io_enq_bits_data_addr_beat;
  wire  roq_io_enq_bits_data_subblock;
  wire [1:0] roq_io_enq_bits_tag;
  wire  roq_io_deq_valid;
  wire [1:0] roq_io_deq_tag;
  wire [2:0] roq_io_deq_data_addr_beat;
  wire  roq_io_deq_data_subblock;
  wire  roq_io_deq_matches;
  wire  get_id_mapper_clk;
  wire  get_id_mapper_reset;
  wire  get_id_mapper_io_req_valid;
  wire  get_id_mapper_io_req_ready;
  wire [1:0] get_id_mapper_io_req_in_id;
  wire [4:0] get_id_mapper_io_req_out_id;
  wire  get_id_mapper_io_resp_valid;
  wire  get_id_mapper_io_resp_matches;
  wire [4:0] get_id_mapper_io_resp_out_id;
  wire [1:0] get_id_mapper_io_resp_in_id;
  wire  put_id_mapper_clk;
  wire  put_id_mapper_reset;
  wire  put_id_mapper_io_req_valid;
  wire  put_id_mapper_io_req_ready;
  wire [1:0] put_id_mapper_io_req_in_id;
  wire [4:0] put_id_mapper_io_req_out_id;
  wire  put_id_mapper_io_resp_valid;
  wire  put_id_mapper_io_resp_matches;
  wire [4:0] put_id_mapper_io_resp_out_id;
  wire [1:0] put_id_mapper_io_resp_in_id;
  wire  T_755;
  wire  put_id_mask;
  wire  T_757;
  wire  put_id_ready;
  reg  w_inflight;
  reg [31:0] GEN_12;
  reg [4:0] w_id_reg;
  reg [31:0] GEN_13;
  wire [4:0] w_id;
  wire  aw_ready;
  wire  T_760;
  wire  T_762;
  wire  T_763;
  reg [2:0] nasti_cnt_out;
  reg [31:0] GEN_14;
  wire  T_766;
  wire [3:0] T_768;
  wire [2:0] T_769;
  wire [2:0] GEN_1;
  wire  nasti_wrap_out;
  wire  T_770;
  wire  T_771;
  wire  T_773;
  wire  T_774;
  wire  T_775;
  wire  T_776;
  wire  T_778;
  wire  T_779;
  wire  T_780;
  wire  T_781;
  wire  T_782;
  wire  T_784;
  wire [2:0] T_792_0;
  wire [2:0] T_792_1;
  wire  T_794;
  wire  T_795;
  wire  T_796;
  wire  T_797;
  wire [2:0] T_798;
  wire [2:0] T_800;
  wire [28:0] T_801;
  wire [31:0] T_802;
  wire [1:0] T_803;
  wire [1:0] T_805;
  wire [2:0] T_808;
  wire [31:0] T_821_addr;
  wire [7:0] T_821_len;
  wire [2:0] T_821_size;
  wire [1:0] T_821_burst;
  wire  T_821_lock;
  wire [3:0] T_821_cache;
  wire [2:0] T_821_prot;
  wire [3:0] T_821_qos;
  wire [3:0] T_821_region;
  wire [4:0] T_821_id;
  wire  T_821_user;
  wire  T_840;
  wire  T_841;
  wire  T_865;
  wire  T_866;
  wire  T_868;
  wire  T_869;
  wire  T_870;
  wire [7:0] T_871;
  wire [7:0] T_873;
  wire [7:0] T_874;
  wire [7:0] T_875;
  wire  all_inside_0_0;
  wire  all_inside_0_1;
  wire  all_inside_0_2;
  wire  all_inside_0_3;
  wire  all_inside_0_4;
  wire  all_inside_0_5;
  wire  all_inside_0_6;
  wire  all_inside_0_7;
  wire  T_876;
  wire  T_877;
  wire  T_878;
  wire  T_879;
  wire  T_880;
  wire  T_881;
  wire  T_888;
  wire [1:0] T_889;
  wire [1:0] T_891;
  wire  T_892;
  wire  T_893;
  wire  T_894;
  wire  T_895;
  wire  T_896;
  wire  T_897;
  wire  T_898;
  wire  T_899;
  wire [2:0] T_900;
  wire [1:0] T_902;
  wire  T_903;
  wire  T_904;
  wire  T_905;
  wire  T_906;
  wire  T_907;
  wire  T_908;
  wire  T_909;
  wire  T_910;
  wire  T_911;
  wire  T_912;
  wire  T_913;
  wire  T_914;
  wire  T_915;
  wire  T_916;
  wire  T_917;
  wire  T_918;
  wire  T_919;
  wire  T_920;
  wire [3:0] put_offset;
  wire [1:0] put_size;
  wire  T_923;
  wire  T_924;
  wire  T_925;
  wire  T_926;
  wire [2:0] T_934_0;
  wire [2:0] T_934_1;
  wire  T_936;
  wire  T_937;
  wire  T_938;
  wire  T_939;
  wire [2:0] T_942;
  wire [31:0] T_944;
  wire [3:0] T_946;
  wire [31:0] GEN_7;
  wire [31:0] T_947;
  wire [1:0] T_949;
  wire [2:0] T_952;
  wire [31:0] T_965_addr;
  wire [7:0] T_965_len;
  wire [2:0] T_965_size;
  wire [1:0] T_965_burst;
  wire  T_965_lock;
  wire [3:0] T_965_cache;
  wire [2:0] T_965_prot;
  wire [3:0] T_965_qos;
  wire [3:0] T_965_region;
  wire [4:0] T_965_id;
  wire  T_965_user;
  wire  T_984;
  wire  T_1024;
  wire  T_1025;
  wire [63:0] T_1032_data;
  wire  T_1032_last;
  wire [4:0] T_1032_id;
  wire [7:0] T_1032_strb;
  wire  T_1032_user;
  wire  T_1039;
  wire  T_1040;
  wire  T_1041;
  wire  T_1042;
  wire  T_1043;
  wire  T_1047;
  wire  T_1048;
  wire  GEN_2;
  wire [4:0] GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  T_1051;
  wire [2:0] T_1059_0;
  wire [3:0] GEN_8;
  wire  T_1061;
  wire  T_1062;
  wire  T_1063;
  wire  T_1065;
  reg [2:0] tl_cnt_in;
  reg [31:0] GEN_15;
  wire [3:0] T_1070;
  wire [2:0] T_1071;
  wire [2:0] GEN_6;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_0_bits_client_id;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_1_bits_client_id;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_out_bits_client_id;
  wire  gnt_arb_io_chosen;
  wire [2:0] T_1103;
  wire [2:0] T_1105;
  wire [2:0] T_1133_addr_beat;
  wire [1:0] T_1133_client_xact_id;
  wire  T_1133_manager_xact_id;
  wire  T_1133_is_builtin_type;
  wire [3:0] T_1133_g_type;
  wire [63:0] T_1133_data;
  wire  T_1161;
  wire  T_1162;
  wire  T_1163;
  wire  T_1165;
  wire  T_1167;
  wire  T_1168;
  wire  T_1169;
  wire  T_1171;
  wire [2:0] T_1204_addr_beat;
  wire [1:0] T_1204_client_xact_id;
  wire  T_1204_manager_xact_id;
  wire  T_1204_is_builtin_type;
  wire [3:0] T_1204_g_type;
  wire [63:0] T_1204_data;
  wire  T_1232;
  wire  T_1233;
  wire  T_1234;
  wire  T_1236;
  wire  T_1238;
  wire  T_1240;
  wire  T_1241;
  wire  T_1242;
  wire  T_1244;
  wire  T_1246;
  wire  T_1248;
  wire  T_1249;
  wire  T_1250;
  wire  T_1252;
  wire  GEN_9;
  reg [31:0] GEN_16;
  wire  GEN_10;
  reg [31:0] GEN_17;
  ReorderQueue_2 roq (
    .clk(roq_clk),
    .reset(roq_reset),
    .io_enq_ready(roq_io_enq_ready),
    .io_enq_valid(roq_io_enq_valid),
    .io_enq_bits_data_addr_beat(roq_io_enq_bits_data_addr_beat),
    .io_enq_bits_data_subblock(roq_io_enq_bits_data_subblock),
    .io_enq_bits_tag(roq_io_enq_bits_tag),
    .io_deq_valid(roq_io_deq_valid),
    .io_deq_tag(roq_io_deq_tag),
    .io_deq_data_addr_beat(roq_io_deq_data_addr_beat),
    .io_deq_data_subblock(roq_io_deq_data_subblock),
    .io_deq_matches(roq_io_deq_matches)
  );
  IdMapper get_id_mapper (
    .clk(get_id_mapper_clk),
    .reset(get_id_mapper_reset),
    .io_req_valid(get_id_mapper_io_req_valid),
    .io_req_ready(get_id_mapper_io_req_ready),
    .io_req_in_id(get_id_mapper_io_req_in_id),
    .io_req_out_id(get_id_mapper_io_req_out_id),
    .io_resp_valid(get_id_mapper_io_resp_valid),
    .io_resp_matches(get_id_mapper_io_resp_matches),
    .io_resp_out_id(get_id_mapper_io_resp_out_id),
    .io_resp_in_id(get_id_mapper_io_resp_in_id)
  );
  IdMapper put_id_mapper (
    .clk(put_id_mapper_clk),
    .reset(put_id_mapper_reset),
    .io_req_valid(put_id_mapper_io_req_valid),
    .io_req_ready(put_id_mapper_io_req_ready),
    .io_req_in_id(put_id_mapper_io_req_in_id),
    .io_req_out_id(put_id_mapper_io_req_out_id),
    .io_resp_valid(put_id_mapper_io_resp_valid),
    .io_resp_matches(put_id_mapper_io_resp_matches),
    .io_resp_out_id(put_id_mapper_io_resp_out_id),
    .io_resp_in_id(put_id_mapper_io_resp_in_id)
  );
  LockingArbiter gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_0_bits_client_id(gnt_arb_io_in_0_bits_client_id),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_1_bits_client_id(gnt_arb_io_in_1_bits_client_id),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_out_bits_client_id(gnt_arb_io_out_bits_client_id),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_tl_acquire_ready = T_1043;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_nasti_aw_valid = T_926;
  assign io_nasti_aw_bits_addr = T_965_addr;
  assign io_nasti_aw_bits_len = T_965_len;
  assign io_nasti_aw_bits_size = T_965_size;
  assign io_nasti_aw_bits_burst = T_965_burst;
  assign io_nasti_aw_bits_lock = T_965_lock;
  assign io_nasti_aw_bits_cache = T_965_cache;
  assign io_nasti_aw_bits_prot = T_965_prot;
  assign io_nasti_aw_bits_qos = T_965_qos;
  assign io_nasti_aw_bits_region = T_965_region;
  assign io_nasti_aw_bits_id = T_965_id;
  assign io_nasti_aw_bits_user = T_965_user;
  assign io_nasti_w_valid = T_984;
  assign io_nasti_w_bits_data = T_1032_data;
  assign io_nasti_w_bits_last = T_1032_last;
  assign io_nasti_w_bits_id = T_1032_id;
  assign io_nasti_w_bits_strb = T_1032_strb;
  assign io_nasti_w_bits_user = T_1032_user;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_ar_valid = T_784;
  assign io_nasti_ar_bits_addr = T_821_addr;
  assign io_nasti_ar_bits_len = T_821_len;
  assign io_nasti_ar_bits_size = T_821_size;
  assign io_nasti_ar_bits_burst = T_821_burst;
  assign io_nasti_ar_bits_lock = T_821_lock;
  assign io_nasti_ar_bits_cache = T_821_cache;
  assign io_nasti_ar_bits_prot = T_821_prot;
  assign io_nasti_ar_bits_qos = T_821_qos;
  assign io_nasti_ar_bits_region = T_821_region;
  assign io_nasti_ar_bits_id = T_821_id;
  assign io_nasti_ar_bits_user = T_821_user;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign T_688_0 = 3'h2;
  assign T_688_1 = 3'h3;
  assign T_688_2 = 3'h4;
  assign T_690 = io_tl_acquire_bits_a_type == T_688_0;
  assign T_691 = io_tl_acquire_bits_a_type == T_688_1;
  assign T_692 = io_tl_acquire_bits_a_type == T_688_2;
  assign T_693 = T_690 | T_691;
  assign T_694 = T_693 | T_692;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T_694;
  assign T_703_0 = 3'h2;
  assign T_703_1 = 3'h0;
  assign T_703_2 = 3'h4;
  assign T_705 = io_tl_acquire_bits_a_type == T_703_0;
  assign T_706 = io_tl_acquire_bits_a_type == T_703_1;
  assign T_707 = io_tl_acquire_bits_a_type == T_703_2;
  assign T_708 = T_705 | T_706;
  assign T_709 = T_708 | T_707;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T_709;
  assign T_718_0 = 3'h3;
  assign T_720 = io_tl_acquire_bits_a_type == T_718_0;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T_720;
  assign T_721 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T_722 = T_721 & is_multibeat;
  assign T_725 = tl_cnt_out == 3'h7;
  assign T_727 = tl_cnt_out + 3'h1;
  assign T_728 = T_727[2:0];
  assign GEN_0 = T_722 ? T_728 : tl_cnt_out;
  assign tl_wrap_out = T_722 & T_725;
  assign T_730 = has_data == 1'h0;
  assign get_valid = io_tl_acquire_valid & T_730;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign roq_clk = clk;
  assign roq_reset = reset;
  assign roq_io_enq_valid = T_771;
  assign roq_io_enq_bits_data_addr_beat = io_tl_acquire_bits_addr_beat;
  assign roq_io_enq_bits_data_subblock = is_subblock;
  assign roq_io_enq_bits_tag = io_nasti_ar_bits_id[1:0];
  assign roq_io_deq_valid = T_774;
  assign roq_io_deq_tag = io_nasti_r_bits_id[1:0];
  assign get_id_mapper_clk = clk;
  assign get_id_mapper_reset = reset;
  assign get_id_mapper_io_req_valid = T_776;
  assign get_id_mapper_io_req_in_id = io_tl_acquire_bits_client_xact_id;
  assign get_id_mapper_io_resp_valid = T_778;
  assign get_id_mapper_io_resp_out_id = io_nasti_r_bits_id;
  assign put_id_mapper_clk = clk;
  assign put_id_mapper_reset = reset;
  assign put_id_mapper_io_req_valid = T_781;
  assign put_id_mapper_io_req_in_id = io_tl_acquire_bits_client_xact_id;
  assign put_id_mapper_io_resp_valid = T_782;
  assign put_id_mapper_io_resp_out_id = io_nasti_b_bits_id;
  assign T_755 = io_tl_acquire_bits_addr_beat == 3'h0;
  assign put_id_mask = is_subblock | T_755;
  assign T_757 = put_id_mask == 1'h0;
  assign put_id_ready = put_id_mapper_io_req_ready | T_757;
  assign w_id = w_inflight ? w_id_reg : put_id_mapper_io_req_out_id;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T_760 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_762 = roq_io_deq_data_subblock == 1'h0;
  assign T_763 = T_760 & T_762;
  assign T_766 = nasti_cnt_out == 3'h7;
  assign T_768 = nasti_cnt_out + 3'h1;
  assign T_769 = T_768[2:0];
  assign GEN_1 = T_763 ? T_769 : nasti_cnt_out;
  assign nasti_wrap_out = T_763 & T_766;
  assign T_770 = get_valid & io_nasti_ar_ready;
  assign T_771 = T_770 & get_id_mapper_io_req_ready;
  assign T_773 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign T_774 = T_760 & T_773;
  assign T_775 = get_valid & roq_io_enq_ready;
  assign T_776 = T_775 & io_nasti_ar_ready;
  assign T_778 = T_760 & io_nasti_r_bits_last;
  assign T_779 = put_valid & aw_ready;
  assign T_780 = T_779 & io_nasti_w_ready;
  assign T_781 = T_780 & put_id_mask;
  assign T_782 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_784 = T_775 & get_id_mapper_io_req_ready;
  assign T_792_0 = 3'h0;
  assign T_792_1 = 3'h4;
  assign T_794 = io_tl_acquire_bits_a_type == T_792_0;
  assign T_795 = io_tl_acquire_bits_a_type == T_792_1;
  assign T_796 = T_794 | T_795;
  assign T_797 = io_tl_acquire_bits_is_builtin_type & T_796;
  assign T_798 = io_tl_acquire_bits_union[10:8];
  assign T_800 = T_797 ? T_798 : 3'h0;
  assign T_801 = {io_tl_acquire_bits_addr_block,io_tl_acquire_bits_addr_beat};
  assign T_802 = {T_801,T_800};
  assign T_803 = io_tl_acquire_bits_union[7:6];
  assign T_805 = is_subblock ? T_803 : 2'h3;
  assign T_808 = is_subblock ? 3'h0 : 3'h7;
  assign T_821_addr = T_802;
  assign T_821_len = {{5'd0}, T_808};
  assign T_821_size = {{1'd0}, T_805};
  assign T_821_burst = 2'h1;
  assign T_821_lock = 1'h0;
  assign T_821_cache = 4'h0;
  assign T_821_prot = 3'h0;
  assign T_821_qos = 4'h0;
  assign T_821_region = 4'h0;
  assign T_821_id = get_id_mapper_io_req_out_id;
  assign T_821_user = 1'h0;
  assign T_840 = io_tl_acquire_bits_a_type == 3'h4;
  assign T_841 = io_tl_acquire_bits_is_builtin_type & T_840;
  assign T_865 = io_tl_acquire_bits_a_type == 3'h3;
  assign T_866 = io_tl_acquire_bits_is_builtin_type & T_865;
  assign T_868 = io_tl_acquire_bits_a_type == 3'h2;
  assign T_869 = io_tl_acquire_bits_is_builtin_type & T_868;
  assign T_870 = T_866 | T_869;
  assign T_871 = io_tl_acquire_bits_union[8:1];
  assign T_873 = T_870 ? T_871 : 8'h0;
  assign T_874 = T_841 ? 8'hff : T_873;
  assign T_875 = ~ T_874;
  assign all_inside_0_0 = T_875[0];
  assign all_inside_0_1 = T_875[1];
  assign all_inside_0_2 = T_875[2];
  assign all_inside_0_3 = T_875[3];
  assign all_inside_0_4 = T_875[4];
  assign all_inside_0_5 = T_875[5];
  assign all_inside_0_6 = T_875[6];
  assign all_inside_0_7 = T_875[7];
  assign T_876 = all_inside_0_0 & all_inside_0_1;
  assign T_877 = all_inside_0_2 & all_inside_0_3;
  assign T_878 = all_inside_0_4 & all_inside_0_5;
  assign T_879 = all_inside_0_6 & all_inside_0_7;
  assign T_880 = T_876 & T_877;
  assign T_881 = T_878 & T_879;
  assign T_888 = T_881 | T_880;
  assign T_889 = {1'h0,T_880};
  assign T_891 = T_888 ? 2'h2 : 2'h3;
  assign T_892 = T_881 & T_877;
  assign T_893 = T_881 & T_876;
  assign T_894 = T_880 & T_879;
  assign T_895 = T_880 & T_878;
  assign T_896 = T_893 | T_895;
  assign T_897 = T_892 | T_893;
  assign T_898 = T_897 | T_894;
  assign T_899 = T_898 | T_895;
  assign T_900 = {T_889,T_896};
  assign T_902 = T_899 ? 2'h1 : T_891;
  assign T_903 = T_892 & all_inside_0_1;
  assign T_904 = T_892 & all_inside_0_0;
  assign T_905 = T_893 & all_inside_0_3;
  assign T_906 = T_893 & all_inside_0_2;
  assign T_907 = T_894 & all_inside_0_5;
  assign T_908 = T_894 & all_inside_0_4;
  assign T_909 = T_895 & all_inside_0_7;
  assign T_910 = T_895 & all_inside_0_6;
  assign T_911 = T_904 | T_906;
  assign T_912 = T_911 | T_908;
  assign T_913 = T_912 | T_910;
  assign T_914 = T_903 | T_904;
  assign T_915 = T_914 | T_905;
  assign T_916 = T_915 | T_906;
  assign T_917 = T_916 | T_907;
  assign T_918 = T_917 | T_908;
  assign T_919 = T_918 | T_909;
  assign T_920 = T_919 | T_910;
  assign put_offset = {T_900,T_913};
  assign put_size = T_920 ? 2'h0 : T_902;
  assign T_923 = w_inflight == 1'h0;
  assign T_924 = put_valid & io_nasti_w_ready;
  assign T_925 = T_924 & put_id_ready;
  assign T_926 = T_925 & T_923;
  assign T_934_0 = 3'h0;
  assign T_934_1 = 3'h4;
  assign T_936 = io_tl_acquire_bits_a_type == T_934_0;
  assign T_937 = io_tl_acquire_bits_a_type == T_934_1;
  assign T_938 = T_936 | T_937;
  assign T_939 = io_tl_acquire_bits_is_builtin_type & T_938;
  assign T_942 = T_939 ? T_798 : 3'h0;
  assign T_944 = {T_801,T_942};
  assign T_946 = is_multibeat ? 4'h0 : put_offset;
  assign GEN_7 = {{28'd0}, T_946};
  assign T_947 = T_944 | GEN_7;
  assign T_949 = is_multibeat ? 2'h3 : put_size;
  assign T_952 = is_multibeat ? 3'h7 : 3'h0;
  assign T_965_addr = T_947;
  assign T_965_len = {{5'd0}, T_952};
  assign T_965_size = {{1'd0}, T_949};
  assign T_965_burst = 2'h1;
  assign T_965_lock = 1'h0;
  assign T_965_cache = 4'h0;
  assign T_965_prot = 3'h0;
  assign T_965_qos = 4'h0;
  assign T_965_region = 4'h0;
  assign T_965_id = put_id_mapper_io_req_out_id;
  assign T_965_user = 1'h0;
  assign T_984 = T_779 & put_id_ready;
  assign T_1024 = is_multibeat == 1'h0;
  assign T_1025 = w_inflight ? T_725 : T_1024;
  assign T_1032_data = io_tl_acquire_bits_data;
  assign T_1032_last = T_1025;
  assign T_1032_id = w_id;
  assign T_1032_strb = T_874;
  assign T_1032_user = 1'h0;
  assign T_1039 = aw_ready & io_nasti_w_ready;
  assign T_1040 = T_1039 & put_id_ready;
  assign T_1041 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T_1042 = T_1041 & get_id_mapper_io_req_ready;
  assign T_1043 = has_data ? T_1040 : T_1042;
  assign T_1047 = T_923 & T_721;
  assign T_1048 = T_1047 & is_multibeat;
  assign GEN_2 = T_1048 ? 1'h1 : w_inflight;
  assign GEN_3 = T_1048 ? w_id : w_id_reg;
  assign GEN_4 = tl_wrap_out ? 1'h0 : GEN_2;
  assign GEN_5 = w_inflight ? GEN_4 : GEN_2;
  assign T_1051 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_1059_0 = 3'h5;
  assign GEN_8 = {{1'd0}, T_1059_0};
  assign T_1061 = io_tl_grant_bits_g_type == GEN_8;
  assign T_1062 = io_tl_grant_bits_g_type == 4'h0;
  assign T_1063 = io_tl_grant_bits_is_builtin_type ? T_1061 : T_1062;
  assign T_1065 = T_1051 & T_1063;
  assign T_1070 = tl_cnt_in + 3'h1;
  assign T_1071 = T_1070[2:0];
  assign GEN_6 = T_1065 ? T_1071 : tl_cnt_in;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_nasti_r_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = T_1133_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = T_1133_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = T_1133_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = T_1133_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = T_1133_g_type;
  assign gnt_arb_io_in_0_bits_data = T_1133_data;
  assign gnt_arb_io_in_0_bits_client_id = GEN_9;
  assign gnt_arb_io_in_1_valid = io_nasti_b_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = T_1204_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = T_1204_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = T_1204_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = T_1204_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = T_1204_g_type;
  assign gnt_arb_io_in_1_bits_data = T_1204_data;
  assign gnt_arb_io_in_1_bits_client_id = GEN_10;
  assign gnt_arb_io_out_ready = io_tl_grant_ready;
  assign T_1103 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T_1105 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T_1133_addr_beat = T_1105;
  assign T_1133_client_xact_id = get_id_mapper_io_resp_in_id;
  assign T_1133_manager_xact_id = 1'h0;
  assign T_1133_is_builtin_type = 1'h1;
  assign T_1133_g_type = {{1'd0}, T_1103};
  assign T_1133_data = io_nasti_r_bits_data;
  assign T_1161 = roq_io_deq_valid == 1'h0;
  assign T_1162 = T_1161 | roq_io_deq_matches;
  assign T_1163 = T_1162 | reset;
  assign T_1165 = T_1163 == 1'h0;
  assign T_1167 = gnt_arb_io_in_0_valid == 1'h0;
  assign T_1168 = T_1167 | get_id_mapper_io_resp_matches;
  assign T_1169 = T_1168 | reset;
  assign T_1171 = T_1169 == 1'h0;
  assign T_1204_addr_beat = 3'h0;
  assign T_1204_client_xact_id = put_id_mapper_io_resp_in_id;
  assign T_1204_manager_xact_id = 1'h0;
  assign T_1204_is_builtin_type = 1'h1;
  assign T_1204_g_type = 4'h3;
  assign T_1204_data = 64'h0;
  assign T_1232 = gnt_arb_io_in_1_valid == 1'h0;
  assign T_1233 = T_1232 | put_id_mapper_io_resp_matches;
  assign T_1234 = T_1233 | reset;
  assign T_1236 = T_1234 == 1'h0;
  assign T_1238 = io_nasti_r_valid == 1'h0;
  assign T_1240 = io_nasti_r_bits_resp == 2'h0;
  assign T_1241 = T_1238 | T_1240;
  assign T_1242 = T_1241 | reset;
  assign T_1244 = T_1242 == 1'h0;
  assign T_1246 = io_nasti_b_valid == 1'h0;
  assign T_1248 = io_nasti_b_bits_resp == 2'h0;
  assign T_1249 = T_1246 | T_1248;
  assign T_1250 = T_1249 | reset;
  assign T_1252 = T_1250 == 1'h0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_9 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_10 = GEN_17[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_11 = {1{$random}};
  tl_cnt_out = GEN_11[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_12 = {1{$random}};
  w_inflight = GEN_12[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_13 = {1{$random}};
  w_id_reg = GEN_13[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_14 = {1{$random}};
  nasti_cnt_out = GEN_14[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_15 = {1{$random}};
  tl_cnt_in = GEN_15[2:0];
  `endif
  GEN_16 = {1{$random}};
  GEN_17 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else begin
      if(T_722) begin
        tl_cnt_out <= T_728;
      end
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else begin
      if(w_inflight) begin
        if(tl_wrap_out) begin
          w_inflight <= 1'h0;
        end else begin
          if(T_1048) begin
            w_inflight <= 1'h1;
          end
        end
      end else begin
        if(T_1048) begin
          w_inflight <= 1'h1;
        end
      end
    end
    if(reset) begin
      w_id_reg <= 5'h0;
    end else begin
      if(T_1048) begin
        if(w_inflight) begin
        end else begin
          w_id_reg <= put_id_mapper_io_req_out_id;
        end
      end
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else begin
      if(T_763) begin
        nasti_cnt_out <= T_769;
      end
    end
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else begin
      if(T_1065) begin
        tl_cnt_in <= T_1071;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1165) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI converter ReorderQueue: NASTI tag error\n    at Nasti.scala:220 assert(!roq.io.deq.valid || roq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1171) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI ID Mapper: NASTI tag error\n    at Nasti.scala:222 assert(!gnt_arb.io.in(0).valid || get_id_mapper.io.resp.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1236) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at Nasti.scala:234 assert(!gnt_arb.io.in(1).valid || put_id_mapper.io.resp.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1244) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI read error\n    at Nasti.scala:236 assert(!io.nasti.r.valid || io.nasti.r.bits.resp === UInt(0), \"NASTI read error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1252) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI write error\n    at Nasti.scala:237 assert(!io.nasti.b.valid || io.nasti.b.bits.resp === UInt(0), \"NASTI write error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_15(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0] io_enq_bits_len,
  input  [2:0] io_enq_bits_size,
  input  [1:0] io_enq_bits_burst,
  input   io_enq_bits_lock,
  input  [3:0] io_enq_bits_cache,
  input  [2:0] io_enq_bits_prot,
  input  [3:0] io_enq_bits_qos,
  input  [3:0] io_enq_bits_region,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [1:0] io_deq_bits_burst,
  output  io_deq_bits_lock,
  output [3:0] io_deq_bits_cache,
  output [2:0] io_deq_bits_prot,
  output [3:0] io_deq_bits_qos,
  output [3:0] io_deq_bits_region,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [31:0] ram_addr [0:0];
  reg [31:0] GEN_0;
  wire [31:0] ram_addr_T_144_data;
  wire  ram_addr_T_144_addr;
  wire  ram_addr_T_144_en;
  wire [31:0] ram_addr_T_125_data;
  wire  ram_addr_T_125_addr;
  wire  ram_addr_T_125_mask;
  wire  ram_addr_T_125_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] GEN_1;
  wire [7:0] ram_len_T_144_data;
  wire  ram_len_T_144_addr;
  wire  ram_len_T_144_en;
  wire [7:0] ram_len_T_125_data;
  wire  ram_len_T_125_addr;
  wire  ram_len_T_125_mask;
  wire  ram_len_T_125_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_size_T_144_data;
  wire  ram_size_T_144_addr;
  wire  ram_size_T_144_en;
  wire [2:0] ram_size_T_125_data;
  wire  ram_size_T_125_addr;
  wire  ram_size_T_125_mask;
  wire  ram_size_T_125_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_burst_T_144_data;
  wire  ram_burst_T_144_addr;
  wire  ram_burst_T_144_en;
  wire [1:0] ram_burst_T_125_data;
  wire  ram_burst_T_125_addr;
  wire  ram_burst_T_125_mask;
  wire  ram_burst_T_125_en;
  reg  ram_lock [0:0];
  reg [31:0] GEN_4;
  wire  ram_lock_T_144_data;
  wire  ram_lock_T_144_addr;
  wire  ram_lock_T_144_en;
  wire  ram_lock_T_125_data;
  wire  ram_lock_T_125_addr;
  wire  ram_lock_T_125_mask;
  wire  ram_lock_T_125_en;
  reg [3:0] ram_cache [0:0];
  reg [31:0] GEN_5;
  wire [3:0] ram_cache_T_144_data;
  wire  ram_cache_T_144_addr;
  wire  ram_cache_T_144_en;
  wire [3:0] ram_cache_T_125_data;
  wire  ram_cache_T_125_addr;
  wire  ram_cache_T_125_mask;
  wire  ram_cache_T_125_en;
  reg [2:0] ram_prot [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_prot_T_144_data;
  wire  ram_prot_T_144_addr;
  wire  ram_prot_T_144_en;
  wire [2:0] ram_prot_T_125_data;
  wire  ram_prot_T_125_addr;
  wire  ram_prot_T_125_mask;
  wire  ram_prot_T_125_en;
  reg [3:0] ram_qos [0:0];
  reg [31:0] GEN_7;
  wire [3:0] ram_qos_T_144_data;
  wire  ram_qos_T_144_addr;
  wire  ram_qos_T_144_en;
  wire [3:0] ram_qos_T_125_data;
  wire  ram_qos_T_125_addr;
  wire  ram_qos_T_125_mask;
  wire  ram_qos_T_125_en;
  reg [3:0] ram_region [0:0];
  reg [31:0] GEN_8;
  wire [3:0] ram_region_T_144_data;
  wire  ram_region_T_144_addr;
  wire  ram_region_T_144_en;
  wire [3:0] ram_region_T_125_data;
  wire  ram_region_T_125_addr;
  wire  ram_region_T_125_mask;
  wire  ram_region_T_125_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_9;
  wire [4:0] ram_id_T_144_data;
  wire  ram_id_T_144_addr;
  wire  ram_id_T_144_en;
  wire [4:0] ram_id_T_125_data;
  wire  ram_id_T_125_addr;
  wire  ram_id_T_125_mask;
  wire  ram_id_T_125_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_10;
  wire  ram_user_T_144_data;
  wire  ram_user_T_144_addr;
  wire  ram_user_T_144_en;
  wire  ram_user_T_125_data;
  wire  ram_user_T_125_addr;
  wire  ram_user_T_125_mask;
  wire  ram_user_T_125_en;
  reg  maybe_full;
  reg [31:0] GEN_11;
  wire  T_122;
  wire  T_123;
  wire  do_enq;
  wire  T_124;
  wire  do_deq;
  wire  T_139;
  wire  GEN_25;
  wire  T_141;
  wire [1:0] T_156;
  wire  ptr_diff;
  wire [1:0] T_158;
  assign io_enq_ready = T_122;
  assign io_deq_valid = T_141;
  assign io_deq_bits_addr = ram_addr_T_144_data;
  assign io_deq_bits_len = ram_len_T_144_data;
  assign io_deq_bits_size = ram_size_T_144_data;
  assign io_deq_bits_burst = ram_burst_T_144_data;
  assign io_deq_bits_lock = ram_lock_T_144_data;
  assign io_deq_bits_cache = ram_cache_T_144_data;
  assign io_deq_bits_prot = ram_prot_T_144_data;
  assign io_deq_bits_qos = ram_qos_T_144_data;
  assign io_deq_bits_region = ram_region_T_144_data;
  assign io_deq_bits_id = ram_id_T_144_data;
  assign io_deq_bits_user = ram_user_T_144_data;
  assign io_count = T_158[0];
  assign ram_addr_T_144_addr = 1'h0;
  assign ram_addr_T_144_en = 1'h1;
  assign ram_addr_T_144_data = ram_addr[ram_addr_T_144_addr];
  assign ram_addr_T_125_data = io_enq_bits_addr;
  assign ram_addr_T_125_addr = 1'h0;
  assign ram_addr_T_125_mask = do_enq;
  assign ram_addr_T_125_en = do_enq;
  assign ram_len_T_144_addr = 1'h0;
  assign ram_len_T_144_en = 1'h1;
  assign ram_len_T_144_data = ram_len[ram_len_T_144_addr];
  assign ram_len_T_125_data = io_enq_bits_len;
  assign ram_len_T_125_addr = 1'h0;
  assign ram_len_T_125_mask = do_enq;
  assign ram_len_T_125_en = do_enq;
  assign ram_size_T_144_addr = 1'h0;
  assign ram_size_T_144_en = 1'h1;
  assign ram_size_T_144_data = ram_size[ram_size_T_144_addr];
  assign ram_size_T_125_data = io_enq_bits_size;
  assign ram_size_T_125_addr = 1'h0;
  assign ram_size_T_125_mask = do_enq;
  assign ram_size_T_125_en = do_enq;
  assign ram_burst_T_144_addr = 1'h0;
  assign ram_burst_T_144_en = 1'h1;
  assign ram_burst_T_144_data = ram_burst[ram_burst_T_144_addr];
  assign ram_burst_T_125_data = io_enq_bits_burst;
  assign ram_burst_T_125_addr = 1'h0;
  assign ram_burst_T_125_mask = do_enq;
  assign ram_burst_T_125_en = do_enq;
  assign ram_lock_T_144_addr = 1'h0;
  assign ram_lock_T_144_en = 1'h1;
  assign ram_lock_T_144_data = ram_lock[ram_lock_T_144_addr];
  assign ram_lock_T_125_data = io_enq_bits_lock;
  assign ram_lock_T_125_addr = 1'h0;
  assign ram_lock_T_125_mask = do_enq;
  assign ram_lock_T_125_en = do_enq;
  assign ram_cache_T_144_addr = 1'h0;
  assign ram_cache_T_144_en = 1'h1;
  assign ram_cache_T_144_data = ram_cache[ram_cache_T_144_addr];
  assign ram_cache_T_125_data = io_enq_bits_cache;
  assign ram_cache_T_125_addr = 1'h0;
  assign ram_cache_T_125_mask = do_enq;
  assign ram_cache_T_125_en = do_enq;
  assign ram_prot_T_144_addr = 1'h0;
  assign ram_prot_T_144_en = 1'h1;
  assign ram_prot_T_144_data = ram_prot[ram_prot_T_144_addr];
  assign ram_prot_T_125_data = io_enq_bits_prot;
  assign ram_prot_T_125_addr = 1'h0;
  assign ram_prot_T_125_mask = do_enq;
  assign ram_prot_T_125_en = do_enq;
  assign ram_qos_T_144_addr = 1'h0;
  assign ram_qos_T_144_en = 1'h1;
  assign ram_qos_T_144_data = ram_qos[ram_qos_T_144_addr];
  assign ram_qos_T_125_data = io_enq_bits_qos;
  assign ram_qos_T_125_addr = 1'h0;
  assign ram_qos_T_125_mask = do_enq;
  assign ram_qos_T_125_en = do_enq;
  assign ram_region_T_144_addr = 1'h0;
  assign ram_region_T_144_en = 1'h1;
  assign ram_region_T_144_data = ram_region[ram_region_T_144_addr];
  assign ram_region_T_125_data = io_enq_bits_region;
  assign ram_region_T_125_addr = 1'h0;
  assign ram_region_T_125_mask = do_enq;
  assign ram_region_T_125_en = do_enq;
  assign ram_id_T_144_addr = 1'h0;
  assign ram_id_T_144_en = 1'h1;
  assign ram_id_T_144_data = ram_id[ram_id_T_144_addr];
  assign ram_id_T_125_data = io_enq_bits_id;
  assign ram_id_T_125_addr = 1'h0;
  assign ram_id_T_125_mask = do_enq;
  assign ram_id_T_125_en = do_enq;
  assign ram_user_T_144_addr = 1'h0;
  assign ram_user_T_144_en = 1'h1;
  assign ram_user_T_144_data = ram_user[ram_user_T_144_addr];
  assign ram_user_T_125_data = io_enq_bits_user;
  assign ram_user_T_125_addr = 1'h0;
  assign ram_user_T_125_mask = do_enq;
  assign ram_user_T_125_en = do_enq;
  assign T_122 = maybe_full == 1'h0;
  assign T_123 = io_enq_ready & io_enq_valid;
  assign do_enq = T_123;
  assign T_124 = io_deq_ready & io_deq_valid;
  assign do_deq = T_124;
  assign T_139 = do_enq != do_deq;
  assign GEN_25 = T_139 ? do_enq : maybe_full;
  assign T_141 = T_122 == 1'h0;
  assign T_156 = 1'h0 - 1'h0;
  assign ptr_diff = T_156[0:0];
  assign T_158 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = GEN_0[31:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = GEN_1[7:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = GEN_3[1:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_lock[initvar] = GEN_4[0:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = GEN_5[3:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = GEN_6[2:0];
  `endif
  GEN_7 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_qos[initvar] = GEN_7[3:0];
  `endif
  GEN_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_region[initvar] = GEN_8[3:0];
  `endif
  GEN_9 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_9[4:0];
  `endif
  GEN_10 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_10[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_11 = {1{$random}};
  maybe_full = GEN_11[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_T_125_en & ram_addr_T_125_mask) begin
      ram_addr[ram_addr_T_125_addr] <= ram_addr_T_125_data;
    end
    if(ram_len_T_125_en & ram_len_T_125_mask) begin
      ram_len[ram_len_T_125_addr] <= ram_len_T_125_data;
    end
    if(ram_size_T_125_en & ram_size_T_125_mask) begin
      ram_size[ram_size_T_125_addr] <= ram_size_T_125_data;
    end
    if(ram_burst_T_125_en & ram_burst_T_125_mask) begin
      ram_burst[ram_burst_T_125_addr] <= ram_burst_T_125_data;
    end
    if(ram_lock_T_125_en & ram_lock_T_125_mask) begin
      ram_lock[ram_lock_T_125_addr] <= ram_lock_T_125_data;
    end
    if(ram_cache_T_125_en & ram_cache_T_125_mask) begin
      ram_cache[ram_cache_T_125_addr] <= ram_cache_T_125_data;
    end
    if(ram_prot_T_125_en & ram_prot_T_125_mask) begin
      ram_prot[ram_prot_T_125_addr] <= ram_prot_T_125_data;
    end
    if(ram_qos_T_125_en & ram_qos_T_125_mask) begin
      ram_qos[ram_qos_T_125_addr] <= ram_qos_T_125_data;
    end
    if(ram_region_T_125_en & ram_region_T_125_mask) begin
      ram_region[ram_region_T_125_addr] <= ram_region_T_125_data;
    end
    if(ram_id_T_125_en & ram_id_T_125_mask) begin
      ram_id[ram_id_T_125_addr] <= ram_id_T_125_data;
    end
    if(ram_user_T_125_en & ram_user_T_125_mask) begin
      ram_user[ram_user_T_125_addr] <= ram_user_T_125_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_17(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input  [7:0] io_enq_bits_strb,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output [7:0] io_deq_bits_strb,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_0;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_1;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_2;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg [7:0] ram_strb [0:1];
  reg [31:0] GEN_3;
  wire [7:0] ram_strb_T_94_data;
  wire  ram_strb_T_94_addr;
  wire  ram_strb_T_94_en;
  wire [7:0] ram_strb_T_73_data;
  wire  ram_strb_T_73_addr;
  wire  ram_strb_T_73_mask;
  wire  ram_strb_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_strb = ram_strb_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_strb_T_94_addr = T_67;
  assign ram_strb_T_94_en = 1'h1;
  assign ram_strb_T_94_data = ram_strb[ram_strb_T_94_addr];
  assign ram_strb_T_73_data = io_enq_bits_strb;
  assign ram_strb_T_73_addr = T_65;
  assign ram_strb_T_73_mask = do_enq;
  assign ram_strb_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_0[63:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_1[0:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_2[4:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_strb[initvar] = GEN_3[7:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_strb_T_73_en & ram_strb_T_73_mask) begin
      ram_strb[ram_strb_T_73_addr] <= ram_strb_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_65 <= T_83;
      end
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_67 <= T_88;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_89) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_18(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [1:0] ram_resp [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_94_data;
  wire  ram_resp_T_94_addr;
  wire  ram_resp_T_94_en;
  wire [1:0] ram_resp_T_73_data;
  wire  ram_resp_T_73_addr;
  wire  ram_resp_T_73_mask;
  wire  ram_resp_T_73_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_1;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_2;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_3;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_resp = ram_resp_T_94_data;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_resp_T_94_addr = T_67;
  assign ram_resp_T_94_en = 1'h1;
  assign ram_resp_T_94_data = ram_resp[ram_resp_T_94_addr];
  assign ram_resp_T_73_data = io_enq_bits_resp;
  assign ram_resp_T_73_addr = T_65;
  assign ram_resp_T_73_mask = do_enq;
  assign ram_resp_T_73_en = do_enq;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_1[63:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_2[0:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_3[4:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_73_en & ram_resp_T_73_mask) begin
      ram_resp[ram_resp_T_73_addr] <= ram_resp_T_73_data;
    end
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_65 <= T_83;
      end
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_67 <= T_88;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_89) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_19(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [1:0] ram_resp [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_64_data;
  wire  ram_resp_T_64_addr;
  wire  ram_resp_T_64_en;
  wire [1:0] ram_resp_T_53_data;
  wire  ram_resp_T_53_addr;
  wire  ram_resp_T_53_mask;
  wire  ram_resp_T_53_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_1;
  wire [4:0] ram_id_T_64_data;
  wire  ram_id_T_64_addr;
  wire  ram_id_T_64_en;
  wire [4:0] ram_id_T_53_data;
  wire  ram_id_T_53_addr;
  wire  ram_id_T_53_mask;
  wire  ram_id_T_53_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_2;
  wire  ram_user_T_64_data;
  wire  ram_user_T_64_addr;
  wire  ram_user_T_64_en;
  wire  ram_user_T_53_data;
  wire  ram_user_T_53_addr;
  wire  ram_user_T_53_mask;
  wire  ram_user_T_53_en;
  reg  maybe_full;
  reg [31:0] GEN_3;
  wire  T_50;
  wire  T_51;
  wire  do_enq;
  wire  T_52;
  wire  do_deq;
  wire  T_59;
  wire  GEN_9;
  wire  T_61;
  wire [1:0] T_68;
  wire  ptr_diff;
  wire [1:0] T_70;
  assign io_enq_ready = T_50;
  assign io_deq_valid = T_61;
  assign io_deq_bits_resp = ram_resp_T_64_data;
  assign io_deq_bits_id = ram_id_T_64_data;
  assign io_deq_bits_user = ram_user_T_64_data;
  assign io_count = T_70[0];
  assign ram_resp_T_64_addr = 1'h0;
  assign ram_resp_T_64_en = 1'h1;
  assign ram_resp_T_64_data = ram_resp[ram_resp_T_64_addr];
  assign ram_resp_T_53_data = io_enq_bits_resp;
  assign ram_resp_T_53_addr = 1'h0;
  assign ram_resp_T_53_mask = do_enq;
  assign ram_resp_T_53_en = do_enq;
  assign ram_id_T_64_addr = 1'h0;
  assign ram_id_T_64_en = 1'h1;
  assign ram_id_T_64_data = ram_id[ram_id_T_64_addr];
  assign ram_id_T_53_data = io_enq_bits_id;
  assign ram_id_T_53_addr = 1'h0;
  assign ram_id_T_53_mask = do_enq;
  assign ram_id_T_53_en = do_enq;
  assign ram_user_T_64_addr = 1'h0;
  assign ram_user_T_64_en = 1'h1;
  assign ram_user_T_64_data = ram_user[ram_user_T_64_addr];
  assign ram_user_T_53_data = io_enq_bits_user;
  assign ram_user_T_53_addr = 1'h0;
  assign ram_user_T_53_mask = do_enq;
  assign ram_user_T_53_en = do_enq;
  assign T_50 = maybe_full == 1'h0;
  assign T_51 = io_enq_ready & io_enq_valid;
  assign do_enq = T_51;
  assign T_52 = io_deq_ready & io_deq_valid;
  assign do_deq = T_52;
  assign T_59 = do_enq != do_deq;
  assign GEN_9 = T_59 ? do_enq : maybe_full;
  assign T_61 = T_50 == 1'h0;
  assign T_68 = 1'h0 - 1'h0;
  assign ptr_diff = T_68[0:0];
  assign T_70 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_1[4:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  maybe_full = GEN_3[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_53_en & ram_resp_T_53_mask) begin
      ram_resp[ram_resp_T_53_addr] <= ram_resp_T_53_data;
    end
    if(ram_id_T_53_en & ram_id_T_53_mask) begin
      ram_id[ram_id_T_53_addr] <= ram_id_T_53_data;
    end
    if(ram_user_T_53_en & ram_user_T_53_mask) begin
      ram_user[ram_user_T_53_addr] <= ram_user_T_53_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_59) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Periphery(
  input   clk,
  input   reset,
  output  io_mem_in_0_acquire_ready,
  input   io_mem_in_0_acquire_valid,
  input  [25:0] io_mem_in_0_acquire_bits_addr_block,
  input  [1:0] io_mem_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_mem_in_0_acquire_bits_addr_beat,
  input   io_mem_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_mem_in_0_acquire_bits_a_type,
  input  [10:0] io_mem_in_0_acquire_bits_union,
  input  [63:0] io_mem_in_0_acquire_bits_data,
  input   io_mem_in_0_grant_ready,
  output  io_mem_in_0_grant_valid,
  output [2:0] io_mem_in_0_grant_bits_addr_beat,
  output [1:0] io_mem_in_0_grant_bits_client_xact_id,
  output  io_mem_in_0_grant_bits_manager_xact_id,
  output  io_mem_in_0_grant_bits_is_builtin_type,
  output [3:0] io_mem_in_0_grant_bits_g_type,
  output [63:0] io_mem_in_0_grant_bits_data,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user
);
  wire  NastiIOTileLinkIOConverter_1_clk;
  wire  NastiIOTileLinkIOConverter_1_reset;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_ready;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_valid;
  wire [25:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type;
  wire [10:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_ready;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_valid;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_valid;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user;
  wire  Queue_15_1_clk;
  wire  Queue_15_1_reset;
  wire  Queue_15_1_io_enq_ready;
  wire  Queue_15_1_io_enq_valid;
  wire [31:0] Queue_15_1_io_enq_bits_addr;
  wire [7:0] Queue_15_1_io_enq_bits_len;
  wire [2:0] Queue_15_1_io_enq_bits_size;
  wire [1:0] Queue_15_1_io_enq_bits_burst;
  wire  Queue_15_1_io_enq_bits_lock;
  wire [3:0] Queue_15_1_io_enq_bits_cache;
  wire [2:0] Queue_15_1_io_enq_bits_prot;
  wire [3:0] Queue_15_1_io_enq_bits_qos;
  wire [3:0] Queue_15_1_io_enq_bits_region;
  wire [4:0] Queue_15_1_io_enq_bits_id;
  wire  Queue_15_1_io_enq_bits_user;
  wire  Queue_15_1_io_deq_ready;
  wire  Queue_15_1_io_deq_valid;
  wire [31:0] Queue_15_1_io_deq_bits_addr;
  wire [7:0] Queue_15_1_io_deq_bits_len;
  wire [2:0] Queue_15_1_io_deq_bits_size;
  wire [1:0] Queue_15_1_io_deq_bits_burst;
  wire  Queue_15_1_io_deq_bits_lock;
  wire [3:0] Queue_15_1_io_deq_bits_cache;
  wire [2:0] Queue_15_1_io_deq_bits_prot;
  wire [3:0] Queue_15_1_io_deq_bits_qos;
  wire [3:0] Queue_15_1_io_deq_bits_region;
  wire [4:0] Queue_15_1_io_deq_bits_id;
  wire  Queue_15_1_io_deq_bits_user;
  wire  Queue_15_1_io_count;
  wire  Queue_16_1_clk;
  wire  Queue_16_1_reset;
  wire  Queue_16_1_io_enq_ready;
  wire  Queue_16_1_io_enq_valid;
  wire [31:0] Queue_16_1_io_enq_bits_addr;
  wire [7:0] Queue_16_1_io_enq_bits_len;
  wire [2:0] Queue_16_1_io_enq_bits_size;
  wire [1:0] Queue_16_1_io_enq_bits_burst;
  wire  Queue_16_1_io_enq_bits_lock;
  wire [3:0] Queue_16_1_io_enq_bits_cache;
  wire [2:0] Queue_16_1_io_enq_bits_prot;
  wire [3:0] Queue_16_1_io_enq_bits_qos;
  wire [3:0] Queue_16_1_io_enq_bits_region;
  wire [4:0] Queue_16_1_io_enq_bits_id;
  wire  Queue_16_1_io_enq_bits_user;
  wire  Queue_16_1_io_deq_ready;
  wire  Queue_16_1_io_deq_valid;
  wire [31:0] Queue_16_1_io_deq_bits_addr;
  wire [7:0] Queue_16_1_io_deq_bits_len;
  wire [2:0] Queue_16_1_io_deq_bits_size;
  wire [1:0] Queue_16_1_io_deq_bits_burst;
  wire  Queue_16_1_io_deq_bits_lock;
  wire [3:0] Queue_16_1_io_deq_bits_cache;
  wire [2:0] Queue_16_1_io_deq_bits_prot;
  wire [3:0] Queue_16_1_io_deq_bits_qos;
  wire [3:0] Queue_16_1_io_deq_bits_region;
  wire [4:0] Queue_16_1_io_deq_bits_id;
  wire  Queue_16_1_io_deq_bits_user;
  wire  Queue_16_1_io_count;
  wire  Queue_17_1_clk;
  wire  Queue_17_1_reset;
  wire  Queue_17_1_io_enq_ready;
  wire  Queue_17_1_io_enq_valid;
  wire [63:0] Queue_17_1_io_enq_bits_data;
  wire  Queue_17_1_io_enq_bits_last;
  wire [4:0] Queue_17_1_io_enq_bits_id;
  wire [7:0] Queue_17_1_io_enq_bits_strb;
  wire  Queue_17_1_io_enq_bits_user;
  wire  Queue_17_1_io_deq_ready;
  wire  Queue_17_1_io_deq_valid;
  wire [63:0] Queue_17_1_io_deq_bits_data;
  wire  Queue_17_1_io_deq_bits_last;
  wire [4:0] Queue_17_1_io_deq_bits_id;
  wire [7:0] Queue_17_1_io_deq_bits_strb;
  wire  Queue_17_1_io_deq_bits_user;
  wire [1:0] Queue_17_1_io_count;
  wire  Queue_18_1_clk;
  wire  Queue_18_1_reset;
  wire  Queue_18_1_io_enq_ready;
  wire  Queue_18_1_io_enq_valid;
  wire [1:0] Queue_18_1_io_enq_bits_resp;
  wire [63:0] Queue_18_1_io_enq_bits_data;
  wire  Queue_18_1_io_enq_bits_last;
  wire [4:0] Queue_18_1_io_enq_bits_id;
  wire  Queue_18_1_io_enq_bits_user;
  wire  Queue_18_1_io_deq_ready;
  wire  Queue_18_1_io_deq_valid;
  wire [1:0] Queue_18_1_io_deq_bits_resp;
  wire [63:0] Queue_18_1_io_deq_bits_data;
  wire  Queue_18_1_io_deq_bits_last;
  wire [4:0] Queue_18_1_io_deq_bits_id;
  wire  Queue_18_1_io_deq_bits_user;
  wire [1:0] Queue_18_1_io_count;
  wire  Queue_19_1_clk;
  wire  Queue_19_1_reset;
  wire  Queue_19_1_io_enq_ready;
  wire  Queue_19_1_io_enq_valid;
  wire [1:0] Queue_19_1_io_enq_bits_resp;
  wire [4:0] Queue_19_1_io_enq_bits_id;
  wire  Queue_19_1_io_enq_bits_user;
  wire  Queue_19_1_io_deq_ready;
  wire  Queue_19_1_io_deq_valid;
  wire [1:0] Queue_19_1_io_deq_bits_resp;
  wire [4:0] Queue_19_1_io_deq_bits_id;
  wire  Queue_19_1_io_deq_bits_user;
  wire  Queue_19_1_io_count;
  NastiIOTileLinkIOConverter NastiIOTileLinkIOConverter_1 (
    .clk(NastiIOTileLinkIOConverter_1_clk),
    .reset(NastiIOTileLinkIOConverter_1_reset),
    .io_tl_acquire_ready(NastiIOTileLinkIOConverter_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(NastiIOTileLinkIOConverter_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(NastiIOTileLinkIOConverter_1_io_tl_grant_ready),
    .io_tl_grant_valid(NastiIOTileLinkIOConverter_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data),
    .io_nasti_aw_ready(NastiIOTileLinkIOConverter_1_io_nasti_aw_ready),
    .io_nasti_aw_valid(NastiIOTileLinkIOConverter_1_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user),
    .io_nasti_w_ready(NastiIOTileLinkIOConverter_1_io_nasti_w_ready),
    .io_nasti_w_valid(NastiIOTileLinkIOConverter_1_io_nasti_w_valid),
    .io_nasti_w_bits_data(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user),
    .io_nasti_b_ready(NastiIOTileLinkIOConverter_1_io_nasti_b_ready),
    .io_nasti_b_valid(NastiIOTileLinkIOConverter_1_io_nasti_b_valid),
    .io_nasti_b_bits_resp(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user),
    .io_nasti_ar_ready(NastiIOTileLinkIOConverter_1_io_nasti_ar_ready),
    .io_nasti_ar_valid(NastiIOTileLinkIOConverter_1_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user),
    .io_nasti_r_ready(NastiIOTileLinkIOConverter_1_io_nasti_r_ready),
    .io_nasti_r_valid(NastiIOTileLinkIOConverter_1_io_nasti_r_valid),
    .io_nasti_r_bits_resp(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user)
  );
  Queue_15 Queue_15_1 (
    .clk(Queue_15_1_clk),
    .reset(Queue_15_1_reset),
    .io_enq_ready(Queue_15_1_io_enq_ready),
    .io_enq_valid(Queue_15_1_io_enq_valid),
    .io_enq_bits_addr(Queue_15_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_15_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_15_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_15_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_15_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_15_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_15_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_15_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_15_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_15_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_15_1_io_enq_bits_user),
    .io_deq_ready(Queue_15_1_io_deq_ready),
    .io_deq_valid(Queue_15_1_io_deq_valid),
    .io_deq_bits_addr(Queue_15_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_15_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_15_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_15_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_15_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_15_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_15_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_15_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_15_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_15_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_15_1_io_deq_bits_user),
    .io_count(Queue_15_1_io_count)
  );
  Queue_15 Queue_16_1 (
    .clk(Queue_16_1_clk),
    .reset(Queue_16_1_reset),
    .io_enq_ready(Queue_16_1_io_enq_ready),
    .io_enq_valid(Queue_16_1_io_enq_valid),
    .io_enq_bits_addr(Queue_16_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_16_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_16_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_16_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_16_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_16_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_16_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_16_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_16_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_16_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_16_1_io_enq_bits_user),
    .io_deq_ready(Queue_16_1_io_deq_ready),
    .io_deq_valid(Queue_16_1_io_deq_valid),
    .io_deq_bits_addr(Queue_16_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_16_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_16_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_16_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_16_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_16_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_16_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_16_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_16_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_16_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_16_1_io_deq_bits_user),
    .io_count(Queue_16_1_io_count)
  );
  Queue_17 Queue_17_1 (
    .clk(Queue_17_1_clk),
    .reset(Queue_17_1_reset),
    .io_enq_ready(Queue_17_1_io_enq_ready),
    .io_enq_valid(Queue_17_1_io_enq_valid),
    .io_enq_bits_data(Queue_17_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_17_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_17_1_io_enq_bits_id),
    .io_enq_bits_strb(Queue_17_1_io_enq_bits_strb),
    .io_enq_bits_user(Queue_17_1_io_enq_bits_user),
    .io_deq_ready(Queue_17_1_io_deq_ready),
    .io_deq_valid(Queue_17_1_io_deq_valid),
    .io_deq_bits_data(Queue_17_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_17_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_17_1_io_deq_bits_id),
    .io_deq_bits_strb(Queue_17_1_io_deq_bits_strb),
    .io_deq_bits_user(Queue_17_1_io_deq_bits_user),
    .io_count(Queue_17_1_io_count)
  );
  Queue_18 Queue_18_1 (
    .clk(Queue_18_1_clk),
    .reset(Queue_18_1_reset),
    .io_enq_ready(Queue_18_1_io_enq_ready),
    .io_enq_valid(Queue_18_1_io_enq_valid),
    .io_enq_bits_resp(Queue_18_1_io_enq_bits_resp),
    .io_enq_bits_data(Queue_18_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_18_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_18_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_18_1_io_enq_bits_user),
    .io_deq_ready(Queue_18_1_io_deq_ready),
    .io_deq_valid(Queue_18_1_io_deq_valid),
    .io_deq_bits_resp(Queue_18_1_io_deq_bits_resp),
    .io_deq_bits_data(Queue_18_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_18_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_18_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_18_1_io_deq_bits_user),
    .io_count(Queue_18_1_io_count)
  );
  Queue_19 Queue_19_1 (
    .clk(Queue_19_1_clk),
    .reset(Queue_19_1_reset),
    .io_enq_ready(Queue_19_1_io_enq_ready),
    .io_enq_valid(Queue_19_1_io_enq_valid),
    .io_enq_bits_resp(Queue_19_1_io_enq_bits_resp),
    .io_enq_bits_id(Queue_19_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_19_1_io_enq_bits_user),
    .io_deq_ready(Queue_19_1_io_deq_ready),
    .io_deq_valid(Queue_19_1_io_deq_valid),
    .io_deq_bits_resp(Queue_19_1_io_deq_bits_resp),
    .io_deq_bits_id(Queue_19_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_19_1_io_deq_bits_user),
    .io_count(Queue_19_1_io_count)
  );
  assign io_mem_in_0_acquire_ready = NastiIOTileLinkIOConverter_1_io_tl_acquire_ready;
  assign io_mem_in_0_grant_valid = NastiIOTileLinkIOConverter_1_io_tl_grant_valid;
  assign io_mem_in_0_grant_bits_addr_beat = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat;
  assign io_mem_in_0_grant_bits_client_xact_id = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id;
  assign io_mem_in_0_grant_bits_manager_xact_id = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id;
  assign io_mem_in_0_grant_bits_is_builtin_type = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type;
  assign io_mem_in_0_grant_bits_g_type = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type;
  assign io_mem_in_0_grant_bits_data = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data;
  assign io_mem_axi_0_aw_valid = Queue_16_1_io_deq_valid;
  assign io_mem_axi_0_aw_bits_addr = Queue_16_1_io_deq_bits_addr;
  assign io_mem_axi_0_aw_bits_len = Queue_16_1_io_deq_bits_len;
  assign io_mem_axi_0_aw_bits_size = Queue_16_1_io_deq_bits_size;
  assign io_mem_axi_0_aw_bits_burst = Queue_16_1_io_deq_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = Queue_16_1_io_deq_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = 4'h3;
  assign io_mem_axi_0_aw_bits_prot = Queue_16_1_io_deq_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = Queue_16_1_io_deq_bits_qos;
  assign io_mem_axi_0_aw_bits_region = Queue_16_1_io_deq_bits_region;
  assign io_mem_axi_0_aw_bits_id = Queue_16_1_io_deq_bits_id;
  assign io_mem_axi_0_aw_bits_user = Queue_16_1_io_deq_bits_user;
  assign io_mem_axi_0_w_valid = Queue_17_1_io_deq_valid;
  assign io_mem_axi_0_w_bits_data = Queue_17_1_io_deq_bits_data;
  assign io_mem_axi_0_w_bits_last = Queue_17_1_io_deq_bits_last;
  assign io_mem_axi_0_w_bits_id = Queue_17_1_io_deq_bits_id;
  assign io_mem_axi_0_w_bits_strb = Queue_17_1_io_deq_bits_strb;
  assign io_mem_axi_0_w_bits_user = Queue_17_1_io_deq_bits_user;
  assign io_mem_axi_0_b_ready = Queue_19_1_io_enq_ready;
  assign io_mem_axi_0_ar_valid = Queue_15_1_io_deq_valid;
  assign io_mem_axi_0_ar_bits_addr = Queue_15_1_io_deq_bits_addr;
  assign io_mem_axi_0_ar_bits_len = Queue_15_1_io_deq_bits_len;
  assign io_mem_axi_0_ar_bits_size = Queue_15_1_io_deq_bits_size;
  assign io_mem_axi_0_ar_bits_burst = Queue_15_1_io_deq_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = Queue_15_1_io_deq_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = 4'h3;
  assign io_mem_axi_0_ar_bits_prot = Queue_15_1_io_deq_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = Queue_15_1_io_deq_bits_qos;
  assign io_mem_axi_0_ar_bits_region = Queue_15_1_io_deq_bits_region;
  assign io_mem_axi_0_ar_bits_id = Queue_15_1_io_deq_bits_id;
  assign io_mem_axi_0_ar_bits_user = Queue_15_1_io_deq_bits_user;
  assign io_mem_axi_0_r_ready = Queue_18_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_clk = clk;
  assign NastiIOTileLinkIOConverter_1_reset = reset;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_valid = io_mem_in_0_acquire_valid;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block = io_mem_in_0_acquire_bits_addr_block;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id = io_mem_in_0_acquire_bits_client_xact_id;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat = io_mem_in_0_acquire_bits_addr_beat;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type = io_mem_in_0_acquire_bits_is_builtin_type;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type = io_mem_in_0_acquire_bits_a_type;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union = io_mem_in_0_acquire_bits_union;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data = io_mem_in_0_acquire_bits_data;
  assign NastiIOTileLinkIOConverter_1_io_tl_grant_ready = io_mem_in_0_grant_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_aw_ready = Queue_16_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_w_ready = Queue_17_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_valid = Queue_19_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp = Queue_19_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id = Queue_19_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user = Queue_19_1_io_deq_bits_user;
  assign NastiIOTileLinkIOConverter_1_io_nasti_ar_ready = Queue_15_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_valid = Queue_18_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp = Queue_18_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data = Queue_18_1_io_deq_bits_data;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last = Queue_18_1_io_deq_bits_last;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id = Queue_18_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user = Queue_18_1_io_deq_bits_user;
  assign Queue_15_1_clk = clk;
  assign Queue_15_1_reset = reset;
  assign Queue_15_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_ar_valid;
  assign Queue_15_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr;
  assign Queue_15_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len;
  assign Queue_15_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size;
  assign Queue_15_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst;
  assign Queue_15_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock;
  assign Queue_15_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache;
  assign Queue_15_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot;
  assign Queue_15_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos;
  assign Queue_15_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region;
  assign Queue_15_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id;
  assign Queue_15_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user;
  assign Queue_15_1_io_deq_ready = io_mem_axi_0_ar_ready;
  assign Queue_16_1_clk = clk;
  assign Queue_16_1_reset = reset;
  assign Queue_16_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_aw_valid;
  assign Queue_16_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr;
  assign Queue_16_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len;
  assign Queue_16_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size;
  assign Queue_16_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst;
  assign Queue_16_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock;
  assign Queue_16_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache;
  assign Queue_16_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot;
  assign Queue_16_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos;
  assign Queue_16_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region;
  assign Queue_16_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id;
  assign Queue_16_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user;
  assign Queue_16_1_io_deq_ready = io_mem_axi_0_aw_ready;
  assign Queue_17_1_clk = clk;
  assign Queue_17_1_reset = reset;
  assign Queue_17_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_w_valid;
  assign Queue_17_1_io_enq_bits_data = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data;
  assign Queue_17_1_io_enq_bits_last = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last;
  assign Queue_17_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id;
  assign Queue_17_1_io_enq_bits_strb = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb;
  assign Queue_17_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user;
  assign Queue_17_1_io_deq_ready = io_mem_axi_0_w_ready;
  assign Queue_18_1_clk = clk;
  assign Queue_18_1_reset = reset;
  assign Queue_18_1_io_enq_valid = io_mem_axi_0_r_valid;
  assign Queue_18_1_io_enq_bits_resp = io_mem_axi_0_r_bits_resp;
  assign Queue_18_1_io_enq_bits_data = io_mem_axi_0_r_bits_data;
  assign Queue_18_1_io_enq_bits_last = io_mem_axi_0_r_bits_last;
  assign Queue_18_1_io_enq_bits_id = io_mem_axi_0_r_bits_id;
  assign Queue_18_1_io_enq_bits_user = io_mem_axi_0_r_bits_user;
  assign Queue_18_1_io_deq_ready = NastiIOTileLinkIOConverter_1_io_nasti_r_ready;
  assign Queue_19_1_clk = clk;
  assign Queue_19_1_reset = reset;
  assign Queue_19_1_io_enq_valid = io_mem_axi_0_b_valid;
  assign Queue_19_1_io_enq_bits_resp = io_mem_axi_0_b_bits_resp;
  assign Queue_19_1_io_enq_bits_id = io_mem_axi_0_b_bits_id;
  assign Queue_19_1_io_enq_bits_user = io_mem_axi_0_b_bits_user;
  assign Queue_19_1_io_deq_ready = NastiIOTileLinkIOConverter_1_io_nasti_b_ready;
endmodule
module Top_1(
  input   clk,
  input   reset,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  input   io_interrupts_0,
  input   io_interrupts_1,
  output  io_debug_req_ready,
  input   io_debug_req_valid,
  input  [4:0] io_debug_req_bits_addr,
  input  [33:0] io_debug_req_bits_data,
  input  [1:0] io_debug_req_bits_op,
  input   io_debug_resp_ready,
  output  io_debug_resp_valid,
  output [33:0] io_debug_resp_bits_data,
  output [1:0] io_debug_resp_bits_resp
);
  wire  coreplex_clk;
  wire  coreplex_reset;
  wire  coreplex_io_mem_0_acquire_ready;
  wire  coreplex_io_mem_0_acquire_valid;
  wire [25:0] coreplex_io_mem_0_acquire_bits_addr_block;
  wire [1:0] coreplex_io_mem_0_acquire_bits_client_xact_id;
  wire [2:0] coreplex_io_mem_0_acquire_bits_addr_beat;
  wire  coreplex_io_mem_0_acquire_bits_is_builtin_type;
  wire [2:0] coreplex_io_mem_0_acquire_bits_a_type;
  wire [10:0] coreplex_io_mem_0_acquire_bits_union;
  wire [63:0] coreplex_io_mem_0_acquire_bits_data;
  wire  coreplex_io_mem_0_grant_ready;
  wire  coreplex_io_mem_0_grant_valid;
  wire [2:0] coreplex_io_mem_0_grant_bits_addr_beat;
  wire [1:0] coreplex_io_mem_0_grant_bits_client_xact_id;
  wire  coreplex_io_mem_0_grant_bits_manager_xact_id;
  wire  coreplex_io_mem_0_grant_bits_is_builtin_type;
  wire [3:0] coreplex_io_mem_0_grant_bits_g_type;
  wire [63:0] coreplex_io_mem_0_grant_bits_data;
  wire  coreplex_io_interrupts_0;
  wire  coreplex_io_interrupts_1;
  wire  coreplex_io_debug_req_ready;
  wire  coreplex_io_debug_req_valid;
  wire [4:0] coreplex_io_debug_req_bits_addr;
  wire [33:0] coreplex_io_debug_req_bits_data;
  wire [1:0] coreplex_io_debug_req_bits_op;
  wire  coreplex_io_debug_resp_ready;
  wire  coreplex_io_debug_resp_valid;
  wire [33:0] coreplex_io_debug_resp_bits_data;
  wire [1:0] coreplex_io_debug_resp_bits_resp;
  wire  coreplex_io_rtcTick;
  wire  periphery_clk;
  wire  periphery_reset;
  wire  periphery_io_mem_in_0_acquire_ready;
  wire  periphery_io_mem_in_0_acquire_valid;
  wire [25:0] periphery_io_mem_in_0_acquire_bits_addr_block;
  wire [1:0] periphery_io_mem_in_0_acquire_bits_client_xact_id;
  wire [2:0] periphery_io_mem_in_0_acquire_bits_addr_beat;
  wire  periphery_io_mem_in_0_acquire_bits_is_builtin_type;
  wire [2:0] periphery_io_mem_in_0_acquire_bits_a_type;
  wire [10:0] periphery_io_mem_in_0_acquire_bits_union;
  wire [63:0] periphery_io_mem_in_0_acquire_bits_data;
  wire  periphery_io_mem_in_0_grant_ready;
  wire  periphery_io_mem_in_0_grant_valid;
  wire [2:0] periphery_io_mem_in_0_grant_bits_addr_beat;
  wire [1:0] periphery_io_mem_in_0_grant_bits_client_xact_id;
  wire  periphery_io_mem_in_0_grant_bits_manager_xact_id;
  wire  periphery_io_mem_in_0_grant_bits_is_builtin_type;
  wire [3:0] periphery_io_mem_in_0_grant_bits_g_type;
  wire [63:0] periphery_io_mem_in_0_grant_bits_data;
  wire  periphery_io_mem_axi_0_aw_ready;
  wire  periphery_io_mem_axi_0_aw_valid;
  wire [31:0] periphery_io_mem_axi_0_aw_bits_addr;
  wire [7:0] periphery_io_mem_axi_0_aw_bits_len;
  wire [2:0] periphery_io_mem_axi_0_aw_bits_size;
  wire [1:0] periphery_io_mem_axi_0_aw_bits_burst;
  wire  periphery_io_mem_axi_0_aw_bits_lock;
  wire [3:0] periphery_io_mem_axi_0_aw_bits_cache;
  wire [2:0] periphery_io_mem_axi_0_aw_bits_prot;
  wire [3:0] periphery_io_mem_axi_0_aw_bits_qos;
  wire [3:0] periphery_io_mem_axi_0_aw_bits_region;
  wire [4:0] periphery_io_mem_axi_0_aw_bits_id;
  wire  periphery_io_mem_axi_0_aw_bits_user;
  wire  periphery_io_mem_axi_0_w_ready;
  wire  periphery_io_mem_axi_0_w_valid;
  wire [63:0] periphery_io_mem_axi_0_w_bits_data;
  wire  periphery_io_mem_axi_0_w_bits_last;
  wire [4:0] periphery_io_mem_axi_0_w_bits_id;
  wire [7:0] periphery_io_mem_axi_0_w_bits_strb;
  wire  periphery_io_mem_axi_0_w_bits_user;
  wire  periphery_io_mem_axi_0_b_ready;
  wire  periphery_io_mem_axi_0_b_valid;
  wire [1:0] periphery_io_mem_axi_0_b_bits_resp;
  wire [4:0] periphery_io_mem_axi_0_b_bits_id;
  wire  periphery_io_mem_axi_0_b_bits_user;
  wire  periphery_io_mem_axi_0_ar_ready;
  wire  periphery_io_mem_axi_0_ar_valid;
  wire [31:0] periphery_io_mem_axi_0_ar_bits_addr;
  wire [7:0] periphery_io_mem_axi_0_ar_bits_len;
  wire [2:0] periphery_io_mem_axi_0_ar_bits_size;
  wire [1:0] periphery_io_mem_axi_0_ar_bits_burst;
  wire  periphery_io_mem_axi_0_ar_bits_lock;
  wire [3:0] periphery_io_mem_axi_0_ar_bits_cache;
  wire [2:0] periphery_io_mem_axi_0_ar_bits_prot;
  wire [3:0] periphery_io_mem_axi_0_ar_bits_qos;
  wire [3:0] periphery_io_mem_axi_0_ar_bits_region;
  wire [4:0] periphery_io_mem_axi_0_ar_bits_id;
  wire  periphery_io_mem_axi_0_ar_bits_user;
  wire  periphery_io_mem_axi_0_r_ready;
  wire  periphery_io_mem_axi_0_r_valid;
  wire [1:0] periphery_io_mem_axi_0_r_bits_resp;
  wire [63:0] periphery_io_mem_axi_0_r_bits_data;
  wire  periphery_io_mem_axi_0_r_bits_last;
  wire [4:0] periphery_io_mem_axi_0_r_bits_id;
  wire  periphery_io_mem_axi_0_r_bits_user;
  reg [6:0] T_3628;
  reg [31:0] GEN_1;
  wire  T_3630;
  wire [7:0] T_3632;
  wire [6:0] T_3633;
  wire [6:0] GEN_0;
  DefaultCoreplex coreplex (
    .clk(coreplex_clk),
    .reset(coreplex_reset),
    .io_mem_0_acquire_ready(coreplex_io_mem_0_acquire_ready),
    .io_mem_0_acquire_valid(coreplex_io_mem_0_acquire_valid),
    .io_mem_0_acquire_bits_addr_block(coreplex_io_mem_0_acquire_bits_addr_block),
    .io_mem_0_acquire_bits_client_xact_id(coreplex_io_mem_0_acquire_bits_client_xact_id),
    .io_mem_0_acquire_bits_addr_beat(coreplex_io_mem_0_acquire_bits_addr_beat),
    .io_mem_0_acquire_bits_is_builtin_type(coreplex_io_mem_0_acquire_bits_is_builtin_type),
    .io_mem_0_acquire_bits_a_type(coreplex_io_mem_0_acquire_bits_a_type),
    .io_mem_0_acquire_bits_union(coreplex_io_mem_0_acquire_bits_union),
    .io_mem_0_acquire_bits_data(coreplex_io_mem_0_acquire_bits_data),
    .io_mem_0_grant_ready(coreplex_io_mem_0_grant_ready),
    .io_mem_0_grant_valid(coreplex_io_mem_0_grant_valid),
    .io_mem_0_grant_bits_addr_beat(coreplex_io_mem_0_grant_bits_addr_beat),
    .io_mem_0_grant_bits_client_xact_id(coreplex_io_mem_0_grant_bits_client_xact_id),
    .io_mem_0_grant_bits_manager_xact_id(coreplex_io_mem_0_grant_bits_manager_xact_id),
    .io_mem_0_grant_bits_is_builtin_type(coreplex_io_mem_0_grant_bits_is_builtin_type),
    .io_mem_0_grant_bits_g_type(coreplex_io_mem_0_grant_bits_g_type),
    .io_mem_0_grant_bits_data(coreplex_io_mem_0_grant_bits_data),
    .io_interrupts_0(coreplex_io_interrupts_0),
    .io_interrupts_1(coreplex_io_interrupts_1),
    .io_debug_req_ready(coreplex_io_debug_req_ready),
    .io_debug_req_valid(coreplex_io_debug_req_valid),
    .io_debug_req_bits_addr(coreplex_io_debug_req_bits_addr),
    .io_debug_req_bits_data(coreplex_io_debug_req_bits_data),
    .io_debug_req_bits_op(coreplex_io_debug_req_bits_op),
    .io_debug_resp_ready(coreplex_io_debug_resp_ready),
    .io_debug_resp_valid(coreplex_io_debug_resp_valid),
    .io_debug_resp_bits_data(coreplex_io_debug_resp_bits_data),
    .io_debug_resp_bits_resp(coreplex_io_debug_resp_bits_resp),
    .io_rtcTick(coreplex_io_rtcTick)
  );
  Periphery periphery (
    .clk(periphery_clk),
    .reset(periphery_reset),
    .io_mem_in_0_acquire_ready(periphery_io_mem_in_0_acquire_ready),
    .io_mem_in_0_acquire_valid(periphery_io_mem_in_0_acquire_valid),
    .io_mem_in_0_acquire_bits_addr_block(periphery_io_mem_in_0_acquire_bits_addr_block),
    .io_mem_in_0_acquire_bits_client_xact_id(periphery_io_mem_in_0_acquire_bits_client_xact_id),
    .io_mem_in_0_acquire_bits_addr_beat(periphery_io_mem_in_0_acquire_bits_addr_beat),
    .io_mem_in_0_acquire_bits_is_builtin_type(periphery_io_mem_in_0_acquire_bits_is_builtin_type),
    .io_mem_in_0_acquire_bits_a_type(periphery_io_mem_in_0_acquire_bits_a_type),
    .io_mem_in_0_acquire_bits_union(periphery_io_mem_in_0_acquire_bits_union),
    .io_mem_in_0_acquire_bits_data(periphery_io_mem_in_0_acquire_bits_data),
    .io_mem_in_0_grant_ready(periphery_io_mem_in_0_grant_ready),
    .io_mem_in_0_grant_valid(periphery_io_mem_in_0_grant_valid),
    .io_mem_in_0_grant_bits_addr_beat(periphery_io_mem_in_0_grant_bits_addr_beat),
    .io_mem_in_0_grant_bits_client_xact_id(periphery_io_mem_in_0_grant_bits_client_xact_id),
    .io_mem_in_0_grant_bits_manager_xact_id(periphery_io_mem_in_0_grant_bits_manager_xact_id),
    .io_mem_in_0_grant_bits_is_builtin_type(periphery_io_mem_in_0_grant_bits_is_builtin_type),
    .io_mem_in_0_grant_bits_g_type(periphery_io_mem_in_0_grant_bits_g_type),
    .io_mem_in_0_grant_bits_data(periphery_io_mem_in_0_grant_bits_data),
    .io_mem_axi_0_aw_ready(periphery_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(periphery_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(periphery_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(periphery_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(periphery_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(periphery_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(periphery_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(periphery_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(periphery_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(periphery_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(periphery_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(periphery_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(periphery_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(periphery_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(periphery_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(periphery_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(periphery_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(periphery_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(periphery_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(periphery_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(periphery_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(periphery_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(periphery_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(periphery_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(periphery_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(periphery_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(periphery_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(periphery_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(periphery_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(periphery_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(periphery_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(periphery_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(periphery_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(periphery_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(periphery_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(periphery_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(periphery_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(periphery_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(periphery_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(periphery_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(periphery_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(periphery_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(periphery_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(periphery_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(periphery_io_mem_axi_0_r_bits_user)
  );
  assign io_mem_axi_0_aw_valid = periphery_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = periphery_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = periphery_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = periphery_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = periphery_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = periphery_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = periphery_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = periphery_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = periphery_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = periphery_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = periphery_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = periphery_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = periphery_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = periphery_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = periphery_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = periphery_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = periphery_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = periphery_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = periphery_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = periphery_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = periphery_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = periphery_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = periphery_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = periphery_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = periphery_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = periphery_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = periphery_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = periphery_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = periphery_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = periphery_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = periphery_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = periphery_io_mem_axi_0_r_ready;
  assign io_debug_req_ready = coreplex_io_debug_req_ready;
  assign io_debug_resp_valid = coreplex_io_debug_resp_valid;
  assign io_debug_resp_bits_data = coreplex_io_debug_resp_bits_data;
  assign io_debug_resp_bits_resp = coreplex_io_debug_resp_bits_resp;
  assign coreplex_clk = clk;
  assign coreplex_reset = reset;
  assign coreplex_io_mem_0_acquire_ready = periphery_io_mem_in_0_acquire_ready;
  assign coreplex_io_mem_0_grant_valid = periphery_io_mem_in_0_grant_valid;
  assign coreplex_io_mem_0_grant_bits_addr_beat = periphery_io_mem_in_0_grant_bits_addr_beat;
  assign coreplex_io_mem_0_grant_bits_client_xact_id = periphery_io_mem_in_0_grant_bits_client_xact_id;
  assign coreplex_io_mem_0_grant_bits_manager_xact_id = periphery_io_mem_in_0_grant_bits_manager_xact_id;
  assign coreplex_io_mem_0_grant_bits_is_builtin_type = periphery_io_mem_in_0_grant_bits_is_builtin_type;
  assign coreplex_io_mem_0_grant_bits_g_type = periphery_io_mem_in_0_grant_bits_g_type;
  assign coreplex_io_mem_0_grant_bits_data = periphery_io_mem_in_0_grant_bits_data;
  assign coreplex_io_interrupts_0 = io_interrupts_0;
  assign coreplex_io_interrupts_1 = io_interrupts_1;
  assign coreplex_io_debug_req_valid = io_debug_req_valid;
  assign coreplex_io_debug_req_bits_addr = io_debug_req_bits_addr;
  assign coreplex_io_debug_req_bits_data = io_debug_req_bits_data;
  assign coreplex_io_debug_req_bits_op = io_debug_req_bits_op;
  assign coreplex_io_debug_resp_ready = io_debug_resp_ready;
  assign coreplex_io_rtcTick = T_3630;
  assign periphery_clk = clk;
  assign periphery_reset = reset;
  assign periphery_io_mem_in_0_acquire_valid = coreplex_io_mem_0_acquire_valid;
  assign periphery_io_mem_in_0_acquire_bits_addr_block = coreplex_io_mem_0_acquire_bits_addr_block;
  assign periphery_io_mem_in_0_acquire_bits_client_xact_id = coreplex_io_mem_0_acquire_bits_client_xact_id;
  assign periphery_io_mem_in_0_acquire_bits_addr_beat = coreplex_io_mem_0_acquire_bits_addr_beat;
  assign periphery_io_mem_in_0_acquire_bits_is_builtin_type = coreplex_io_mem_0_acquire_bits_is_builtin_type;
  assign periphery_io_mem_in_0_acquire_bits_a_type = coreplex_io_mem_0_acquire_bits_a_type;
  assign periphery_io_mem_in_0_acquire_bits_union = coreplex_io_mem_0_acquire_bits_union;
  assign periphery_io_mem_in_0_acquire_bits_data = coreplex_io_mem_0_acquire_bits_data;
  assign periphery_io_mem_in_0_grant_ready = coreplex_io_mem_0_grant_ready;
  assign periphery_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign periphery_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign periphery_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign periphery_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign periphery_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign periphery_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign periphery_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign periphery_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign periphery_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign periphery_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign periphery_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign periphery_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign periphery_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign T_3630 = T_3628 == 7'h63;
  assign T_3632 = T_3628 + 7'h1;
  assign T_3633 = T_3632[6:0];
  assign GEN_0 = T_3630 ? 7'h0 : T_3633;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_3628 = GEN_1[6:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_3628 <= 7'h0;
    end else begin
      if(T_3630) begin
        T_3628 <= 7'h0;
      end else begin
        T_3628 <= T_3633;
      end
    end
  end
endmodule
module Top(
  input   clk,
  input   reset,
  output  io_ps_axi_slave_aw_ready,
  input   io_ps_axi_slave_aw_valid,
  input  [31:0] io_ps_axi_slave_aw_bits_addr,
  input  [7:0] io_ps_axi_slave_aw_bits_len,
  input  [2:0] io_ps_axi_slave_aw_bits_size,
  input  [1:0] io_ps_axi_slave_aw_bits_burst,
  input   io_ps_axi_slave_aw_bits_lock,
  input  [3:0] io_ps_axi_slave_aw_bits_cache,
  input  [2:0] io_ps_axi_slave_aw_bits_prot,
  input  [3:0] io_ps_axi_slave_aw_bits_qos,
  input  [3:0] io_ps_axi_slave_aw_bits_region,
  input  [11:0] io_ps_axi_slave_aw_bits_id,
  input   io_ps_axi_slave_aw_bits_user,
  output  io_ps_axi_slave_w_ready,
  input   io_ps_axi_slave_w_valid,
  input  [31:0] io_ps_axi_slave_w_bits_data,
  input   io_ps_axi_slave_w_bits_last,
  input  [11:0] io_ps_axi_slave_w_bits_id,
  input  [3:0] io_ps_axi_slave_w_bits_strb,
  input   io_ps_axi_slave_w_bits_user,
  input   io_ps_axi_slave_b_ready,
  output  io_ps_axi_slave_b_valid,
  output [1:0] io_ps_axi_slave_b_bits_resp,
  output [11:0] io_ps_axi_slave_b_bits_id,
  output  io_ps_axi_slave_b_bits_user,
  output  io_ps_axi_slave_ar_ready,
  input   io_ps_axi_slave_ar_valid,
  input  [31:0] io_ps_axi_slave_ar_bits_addr,
  input  [7:0] io_ps_axi_slave_ar_bits_len,
  input  [2:0] io_ps_axi_slave_ar_bits_size,
  input  [1:0] io_ps_axi_slave_ar_bits_burst,
  input   io_ps_axi_slave_ar_bits_lock,
  input  [3:0] io_ps_axi_slave_ar_bits_cache,
  input  [2:0] io_ps_axi_slave_ar_bits_prot,
  input  [3:0] io_ps_axi_slave_ar_bits_qos,
  input  [3:0] io_ps_axi_slave_ar_bits_region,
  input  [11:0] io_ps_axi_slave_ar_bits_id,
  input   io_ps_axi_slave_ar_bits_user,
  input   io_ps_axi_slave_r_ready,
  output  io_ps_axi_slave_r_valid,
  output [1:0] io_ps_axi_slave_r_bits_resp,
  output [31:0] io_ps_axi_slave_r_bits_data,
  output  io_ps_axi_slave_r_bits_last,
  output [11:0] io_ps_axi_slave_r_bits_id,
  output  io_ps_axi_slave_r_bits_user,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user
);
  wire  adapter_clk;
  wire  adapter_reset;
  wire  adapter_io_nasti_aw_ready;
  wire  adapter_io_nasti_aw_valid;
  wire [31:0] adapter_io_nasti_aw_bits_addr;
  wire [7:0] adapter_io_nasti_aw_bits_len;
  wire [2:0] adapter_io_nasti_aw_bits_size;
  wire [1:0] adapter_io_nasti_aw_bits_burst;
  wire  adapter_io_nasti_aw_bits_lock;
  wire [3:0] adapter_io_nasti_aw_bits_cache;
  wire [2:0] adapter_io_nasti_aw_bits_prot;
  wire [3:0] adapter_io_nasti_aw_bits_qos;
  wire [3:0] adapter_io_nasti_aw_bits_region;
  wire [11:0] adapter_io_nasti_aw_bits_id;
  wire  adapter_io_nasti_aw_bits_user;
  wire  adapter_io_nasti_w_ready;
  wire  adapter_io_nasti_w_valid;
  wire [31:0] adapter_io_nasti_w_bits_data;
  wire  adapter_io_nasti_w_bits_last;
  wire [11:0] adapter_io_nasti_w_bits_id;
  wire [3:0] adapter_io_nasti_w_bits_strb;
  wire  adapter_io_nasti_w_bits_user;
  wire  adapter_io_nasti_b_ready;
  wire  adapter_io_nasti_b_valid;
  wire [1:0] adapter_io_nasti_b_bits_resp;
  wire [11:0] adapter_io_nasti_b_bits_id;
  wire  adapter_io_nasti_b_bits_user;
  wire  adapter_io_nasti_ar_ready;
  wire  adapter_io_nasti_ar_valid;
  wire [31:0] adapter_io_nasti_ar_bits_addr;
  wire [7:0] adapter_io_nasti_ar_bits_len;
  wire [2:0] adapter_io_nasti_ar_bits_size;
  wire [1:0] adapter_io_nasti_ar_bits_burst;
  wire  adapter_io_nasti_ar_bits_lock;
  wire [3:0] adapter_io_nasti_ar_bits_cache;
  wire [2:0] adapter_io_nasti_ar_bits_prot;
  wire [3:0] adapter_io_nasti_ar_bits_qos;
  wire [3:0] adapter_io_nasti_ar_bits_region;
  wire [11:0] adapter_io_nasti_ar_bits_id;
  wire  adapter_io_nasti_ar_bits_user;
  wire  adapter_io_nasti_r_ready;
  wire  adapter_io_nasti_r_valid;
  wire [1:0] adapter_io_nasti_r_bits_resp;
  wire [31:0] adapter_io_nasti_r_bits_data;
  wire  adapter_io_nasti_r_bits_last;
  wire [11:0] adapter_io_nasti_r_bits_id;
  wire  adapter_io_nasti_r_bits_user;
  wire  adapter_io_reset;
  wire  adapter_io_debug_req_ready;
  wire  adapter_io_debug_req_valid;
  wire [4:0] adapter_io_debug_req_bits_addr;
  wire [33:0] adapter_io_debug_req_bits_data;
  wire [1:0] adapter_io_debug_req_bits_op;
  wire  adapter_io_debug_resp_ready;
  wire  adapter_io_debug_resp_valid;
  wire [33:0] adapter_io_debug_resp_bits_data;
  wire [1:0] adapter_io_debug_resp_bits_resp;
  wire  rocket_clk;
  wire  rocket_reset;
  wire  rocket_io_mem_axi_0_aw_ready;
  wire  rocket_io_mem_axi_0_aw_valid;
  wire [31:0] rocket_io_mem_axi_0_aw_bits_addr;
  wire [7:0] rocket_io_mem_axi_0_aw_bits_len;
  wire [2:0] rocket_io_mem_axi_0_aw_bits_size;
  wire [1:0] rocket_io_mem_axi_0_aw_bits_burst;
  wire  rocket_io_mem_axi_0_aw_bits_lock;
  wire [3:0] rocket_io_mem_axi_0_aw_bits_cache;
  wire [2:0] rocket_io_mem_axi_0_aw_bits_prot;
  wire [3:0] rocket_io_mem_axi_0_aw_bits_qos;
  wire [3:0] rocket_io_mem_axi_0_aw_bits_region;
  wire [4:0] rocket_io_mem_axi_0_aw_bits_id;
  wire  rocket_io_mem_axi_0_aw_bits_user;
  wire  rocket_io_mem_axi_0_w_ready;
  wire  rocket_io_mem_axi_0_w_valid;
  wire [63:0] rocket_io_mem_axi_0_w_bits_data;
  wire  rocket_io_mem_axi_0_w_bits_last;
  wire [4:0] rocket_io_mem_axi_0_w_bits_id;
  wire [7:0] rocket_io_mem_axi_0_w_bits_strb;
  wire  rocket_io_mem_axi_0_w_bits_user;
  wire  rocket_io_mem_axi_0_b_ready;
  wire  rocket_io_mem_axi_0_b_valid;
  wire [1:0] rocket_io_mem_axi_0_b_bits_resp;
  wire [4:0] rocket_io_mem_axi_0_b_bits_id;
  wire  rocket_io_mem_axi_0_b_bits_user;
  wire  rocket_io_mem_axi_0_ar_ready;
  wire  rocket_io_mem_axi_0_ar_valid;
  wire [31:0] rocket_io_mem_axi_0_ar_bits_addr;
  wire [7:0] rocket_io_mem_axi_0_ar_bits_len;
  wire [2:0] rocket_io_mem_axi_0_ar_bits_size;
  wire [1:0] rocket_io_mem_axi_0_ar_bits_burst;
  wire  rocket_io_mem_axi_0_ar_bits_lock;
  wire [3:0] rocket_io_mem_axi_0_ar_bits_cache;
  wire [2:0] rocket_io_mem_axi_0_ar_bits_prot;
  wire [3:0] rocket_io_mem_axi_0_ar_bits_qos;
  wire [3:0] rocket_io_mem_axi_0_ar_bits_region;
  wire [4:0] rocket_io_mem_axi_0_ar_bits_id;
  wire  rocket_io_mem_axi_0_ar_bits_user;
  wire  rocket_io_mem_axi_0_r_ready;
  wire  rocket_io_mem_axi_0_r_valid;
  wire [1:0] rocket_io_mem_axi_0_r_bits_resp;
  wire [63:0] rocket_io_mem_axi_0_r_bits_data;
  wire  rocket_io_mem_axi_0_r_bits_last;
  wire [4:0] rocket_io_mem_axi_0_r_bits_id;
  wire  rocket_io_mem_axi_0_r_bits_user;
  wire  rocket_io_interrupts_0;
  wire  rocket_io_interrupts_1;
  wire  rocket_io_debug_req_ready;
  wire  rocket_io_debug_req_valid;
  wire [4:0] rocket_io_debug_req_bits_addr;
  wire [33:0] rocket_io_debug_req_bits_data;
  wire [1:0] rocket_io_debug_req_bits_op;
  wire  rocket_io_debug_resp_ready;
  wire  rocket_io_debug_resp_valid;
  wire [33:0] rocket_io_debug_resp_bits_data;
  wire [1:0] rocket_io_debug_resp_bits_resp;
  ZynqAdapter adapter (
    .clk(adapter_clk),
    .reset(adapter_reset),
    .io_nasti_aw_ready(adapter_io_nasti_aw_ready),
    .io_nasti_aw_valid(adapter_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(adapter_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(adapter_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(adapter_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(adapter_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(adapter_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(adapter_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(adapter_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(adapter_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(adapter_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(adapter_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(adapter_io_nasti_aw_bits_user),
    .io_nasti_w_ready(adapter_io_nasti_w_ready),
    .io_nasti_w_valid(adapter_io_nasti_w_valid),
    .io_nasti_w_bits_data(adapter_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(adapter_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(adapter_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(adapter_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(adapter_io_nasti_w_bits_user),
    .io_nasti_b_ready(adapter_io_nasti_b_ready),
    .io_nasti_b_valid(adapter_io_nasti_b_valid),
    .io_nasti_b_bits_resp(adapter_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(adapter_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(adapter_io_nasti_b_bits_user),
    .io_nasti_ar_ready(adapter_io_nasti_ar_ready),
    .io_nasti_ar_valid(adapter_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(adapter_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(adapter_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(adapter_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(adapter_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(adapter_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(adapter_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(adapter_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(adapter_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(adapter_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(adapter_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(adapter_io_nasti_ar_bits_user),
    .io_nasti_r_ready(adapter_io_nasti_r_ready),
    .io_nasti_r_valid(adapter_io_nasti_r_valid),
    .io_nasti_r_bits_resp(adapter_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(adapter_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(adapter_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(adapter_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(adapter_io_nasti_r_bits_user),
    .io_reset(adapter_io_reset),
    .io_debug_req_ready(adapter_io_debug_req_ready),
    .io_debug_req_valid(adapter_io_debug_req_valid),
    .io_debug_req_bits_addr(adapter_io_debug_req_bits_addr),
    .io_debug_req_bits_data(adapter_io_debug_req_bits_data),
    .io_debug_req_bits_op(adapter_io_debug_req_bits_op),
    .io_debug_resp_ready(adapter_io_debug_resp_ready),
    .io_debug_resp_valid(adapter_io_debug_resp_valid),
    .io_debug_resp_bits_data(adapter_io_debug_resp_bits_data),
    .io_debug_resp_bits_resp(adapter_io_debug_resp_bits_resp)
  );
  Top_1 rocket (
    .clk(rocket_clk),
    .reset(rocket_reset),
    .io_mem_axi_0_aw_ready(rocket_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(rocket_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(rocket_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(rocket_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(rocket_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(rocket_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(rocket_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(rocket_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(rocket_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(rocket_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(rocket_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(rocket_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(rocket_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(rocket_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(rocket_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(rocket_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(rocket_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(rocket_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(rocket_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(rocket_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(rocket_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(rocket_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(rocket_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(rocket_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(rocket_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(rocket_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(rocket_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(rocket_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(rocket_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(rocket_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(rocket_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(rocket_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(rocket_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(rocket_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(rocket_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(rocket_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(rocket_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(rocket_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(rocket_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(rocket_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(rocket_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(rocket_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(rocket_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(rocket_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(rocket_io_mem_axi_0_r_bits_user),
    .io_interrupts_0(rocket_io_interrupts_0),
    .io_interrupts_1(rocket_io_interrupts_1),
    .io_debug_req_ready(rocket_io_debug_req_ready),
    .io_debug_req_valid(rocket_io_debug_req_valid),
    .io_debug_req_bits_addr(rocket_io_debug_req_bits_addr),
    .io_debug_req_bits_data(rocket_io_debug_req_bits_data),
    .io_debug_req_bits_op(rocket_io_debug_req_bits_op),
    .io_debug_resp_ready(rocket_io_debug_resp_ready),
    .io_debug_resp_valid(rocket_io_debug_resp_valid),
    .io_debug_resp_bits_data(rocket_io_debug_resp_bits_data),
    .io_debug_resp_bits_resp(rocket_io_debug_resp_bits_resp)
  );
  assign io_ps_axi_slave_aw_ready = adapter_io_nasti_aw_ready;
  assign io_ps_axi_slave_w_ready = adapter_io_nasti_w_ready;
  assign io_ps_axi_slave_b_valid = adapter_io_nasti_b_valid;
  assign io_ps_axi_slave_b_bits_resp = adapter_io_nasti_b_bits_resp;
  assign io_ps_axi_slave_b_bits_id = adapter_io_nasti_b_bits_id;
  assign io_ps_axi_slave_b_bits_user = adapter_io_nasti_b_bits_user;
  assign io_ps_axi_slave_ar_ready = adapter_io_nasti_ar_ready;
  assign io_ps_axi_slave_r_valid = adapter_io_nasti_r_valid;
  assign io_ps_axi_slave_r_bits_resp = adapter_io_nasti_r_bits_resp;
  assign io_ps_axi_slave_r_bits_data = adapter_io_nasti_r_bits_data;
  assign io_ps_axi_slave_r_bits_last = adapter_io_nasti_r_bits_last;
  assign io_ps_axi_slave_r_bits_id = adapter_io_nasti_r_bits_id;
  assign io_ps_axi_slave_r_bits_user = adapter_io_nasti_r_bits_user;
  assign io_mem_axi_0_aw_valid = rocket_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = rocket_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = rocket_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = rocket_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = rocket_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = rocket_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = rocket_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = rocket_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = rocket_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = rocket_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = rocket_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = rocket_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = rocket_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = rocket_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = rocket_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = rocket_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = rocket_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = rocket_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = rocket_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = rocket_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = rocket_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = rocket_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = rocket_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = rocket_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = rocket_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = rocket_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = rocket_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = rocket_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = rocket_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = rocket_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = rocket_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = rocket_io_mem_axi_0_r_ready;
  assign adapter_clk = clk;
  assign adapter_reset = reset;
  assign adapter_io_nasti_aw_valid = io_ps_axi_slave_aw_valid;
  assign adapter_io_nasti_aw_bits_addr = io_ps_axi_slave_aw_bits_addr;
  assign adapter_io_nasti_aw_bits_len = io_ps_axi_slave_aw_bits_len;
  assign adapter_io_nasti_aw_bits_size = io_ps_axi_slave_aw_bits_size;
  assign adapter_io_nasti_aw_bits_burst = io_ps_axi_slave_aw_bits_burst;
  assign adapter_io_nasti_aw_bits_lock = io_ps_axi_slave_aw_bits_lock;
  assign adapter_io_nasti_aw_bits_cache = io_ps_axi_slave_aw_bits_cache;
  assign adapter_io_nasti_aw_bits_prot = io_ps_axi_slave_aw_bits_prot;
  assign adapter_io_nasti_aw_bits_qos = io_ps_axi_slave_aw_bits_qos;
  assign adapter_io_nasti_aw_bits_region = io_ps_axi_slave_aw_bits_region;
  assign adapter_io_nasti_aw_bits_id = io_ps_axi_slave_aw_bits_id;
  assign adapter_io_nasti_aw_bits_user = io_ps_axi_slave_aw_bits_user;
  assign adapter_io_nasti_w_valid = io_ps_axi_slave_w_valid;
  assign adapter_io_nasti_w_bits_data = io_ps_axi_slave_w_bits_data;
  assign adapter_io_nasti_w_bits_last = io_ps_axi_slave_w_bits_last;
  assign adapter_io_nasti_w_bits_id = io_ps_axi_slave_w_bits_id;
  assign adapter_io_nasti_w_bits_strb = io_ps_axi_slave_w_bits_strb;
  assign adapter_io_nasti_w_bits_user = io_ps_axi_slave_w_bits_user;
  assign adapter_io_nasti_b_ready = io_ps_axi_slave_b_ready;
  assign adapter_io_nasti_ar_valid = io_ps_axi_slave_ar_valid;
  assign adapter_io_nasti_ar_bits_addr = io_ps_axi_slave_ar_bits_addr;
  assign adapter_io_nasti_ar_bits_len = io_ps_axi_slave_ar_bits_len;
  assign adapter_io_nasti_ar_bits_size = io_ps_axi_slave_ar_bits_size;
  assign adapter_io_nasti_ar_bits_burst = io_ps_axi_slave_ar_bits_burst;
  assign adapter_io_nasti_ar_bits_lock = io_ps_axi_slave_ar_bits_lock;
  assign adapter_io_nasti_ar_bits_cache = io_ps_axi_slave_ar_bits_cache;
  assign adapter_io_nasti_ar_bits_prot = io_ps_axi_slave_ar_bits_prot;
  assign adapter_io_nasti_ar_bits_qos = io_ps_axi_slave_ar_bits_qos;
  assign adapter_io_nasti_ar_bits_region = io_ps_axi_slave_ar_bits_region;
  assign adapter_io_nasti_ar_bits_id = io_ps_axi_slave_ar_bits_id;
  assign adapter_io_nasti_ar_bits_user = io_ps_axi_slave_ar_bits_user;
  assign adapter_io_nasti_r_ready = io_ps_axi_slave_r_ready;
  assign adapter_io_debug_req_ready = rocket_io_debug_req_ready;
  assign adapter_io_debug_resp_valid = rocket_io_debug_resp_valid;
  assign adapter_io_debug_resp_bits_data = rocket_io_debug_resp_bits_data;
  assign adapter_io_debug_resp_bits_resp = rocket_io_debug_resp_bits_resp;
  assign rocket_clk = clk;
  assign rocket_reset = adapter_io_reset;
  assign rocket_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign rocket_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign rocket_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign rocket_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign rocket_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign rocket_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign rocket_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign rocket_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign rocket_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign rocket_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign rocket_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign rocket_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign rocket_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign rocket_io_interrupts_0 = 1'h0;
  assign rocket_io_interrupts_1 = 1'h0;
  assign rocket_io_debug_req_valid = adapter_io_debug_req_valid;
  assign rocket_io_debug_req_bits_addr = adapter_io_debug_req_bits_addr;
  assign rocket_io_debug_req_bits_data = adapter_io_debug_req_bits_data;
  assign rocket_io_debug_req_bits_op = adapter_io_debug_req_bits_op;
  assign rocket_io_debug_resp_ready = adapter_io_debug_resp_ready;
endmodule
