module BTB(input clk, input reset,
    input [42:0] io_req,
    output io_resp_valid,
    output io_resp_bits_taken,
    output[42:0] io_resp_bits_target,
    output[2:0] io_resp_bits_entry,
    output[3:0] io_resp_bits_bht_index,
    output[1:0] io_resp_bits_bht_value,
    input  io_update_valid,
    input  io_update_bits_prediction_valid,
    input  io_update_bits_prediction_bits_taken,
    input [42:0] io_update_bits_prediction_bits_target,
    input [2:0] io_update_bits_prediction_bits_entry,
    input [3:0] io_update_bits_prediction_bits_bht_index,
    input [1:0] io_update_bits_prediction_bits_bht_value,
    input [42:0] io_update_bits_pc,
    input [42:0] io_update_bits_target,
    input [42:0] io_update_bits_returnAddr,
    input  io_update_bits_taken,
    input  io_update_bits_isJump,
    input  io_update_bits_isCall,
    input  io_update_bits_isReturn,
    input  io_update_bits_incorrectTarget,
    input  io_invalidate
);

  reg[0:0] T0 = 1'b0;
  wire T1;
  wire T2;
  wire T3;
  reg [42:0] R4;
  wire[42:0] T5;
  wire T6;
  wire T7;
  wire updateTarget;
  reg  R8;
  wire T9;
  wire updateValid;
  reg  updateHit;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  reg  R15;
  wire T406;
  wire[1:0] T16;
  wire[1:0] T17;
  reg [1:0] T18 [15:0];
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg [1:0] R25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  reg  R31;
  wire T32;
  wire T33;
  wire T34;
  reg  R35;
  wire T36;
  wire T37;
  reg [3:0] R38;
  wire[3:0] T39;
  wire[3:0] T40;
  wire[3:0] T41;
  reg [3:0] R42;
  wire[3:0] T43;
  wire[3:0] T44;
  wire[2:0] T45;
  wire[3:0] T46;
  wire[2:0] T407;
  wire[1:0] T408;
  wire T409;
  wire[1:0] T410;
  wire[1:0] T411;
  wire[3:0] T412;
  wire[3:0] T413;
  wire[7:0] hits;
  wire[7:0] T48;
  wire[7:0] T49;
  wire[3:0] T50;
  wire[1:0] T51;
  wire T52;
  wire[3:0] T53;
  wire[3:0] pageHit;
  reg [3:0] pageValid;
  wire[3:0] T414;
  wire[3:0] T54;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] pageReplEn;
  wire[3:0] tgtPageReplEn;
  wire[3:0] tgtPageRepl;
  wire[3:0] T57;
  wire[3:0] T415;
  wire T58;
  wire[3:0] T59;
  wire[2:0] T60;
  wire[3:0] idxPageUpdateOH;
  wire[3:0] idxPageRepl;
  wire[3:0] T61;
  reg [1:0] R62;
  wire[1:0] T416;
  wire[1:0] T63;
  wire[1:0] T64;
  wire T65;
  wire doPageRepl;
  wire doIdxPageRepl;
  wire T66;
  wire[3:0] updatePageHit;
  wire[3:0] T67;
  wire[3:0] T68;
  wire[1:0] T69;
  wire T70;
  wire[29:0] T71;
  reg [42:0] R72;
  wire[42:0] T73;
  wire[29:0] T74;
  reg [29:0] pages [3:0];
  wire[29:0] T75;
  wire[29:0] T76;
  wire[29:0] T77;
  wire[29:0] T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire[29:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[29:0] T89;
  wire[29:0] T90;
  wire[29:0] T91;
  wire[29:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire[29:0] T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[29:0] T102;
  wire[1:0] T103;
  wire T104;
  wire[29:0] T105;
  wire T106;
  wire[29:0] T107;
  wire useUpdatePageHit;
  wire samePage;
  wire[29:0] T108;
  wire[29:0] T109;
  wire doTgtPageRepl;
  wire T110;
  wire usePageHit;
  wire[3:0] T111;
  wire[3:0] T112;
  wire T113;
  wire T114;
  wire[3:0] idxPageReplEn;
  wire T115;
  wire[3:0] T116;
  wire[3:0] T117;
  wire[1:0] T118;
  wire T119;
  wire[29:0] T120;
  wire[29:0] T121;
  wire T122;
  wire[29:0] T123;
  wire[1:0] T124;
  wire T125;
  wire[29:0] T126;
  wire T127;
  wire[29:0] T128;
  wire[3:0] idxPagesOH_0;
  wire[3:0] T129;
  wire[1:0] T130;
  reg [1:0] idxPages [7:0];
  wire[1:0] T131;
  wire[1:0] T417;
  wire T418;
  wire[1:0] T419;
  wire[1:0] T420;
  wire[1:0] T421;
  wire T422;
  wire[2:0] T132;
  reg [2:0] R133;
  wire[2:0] T423;
  wire[2:0] T134;
  wire[2:0] T135;
  wire T136;
  wire T137;
  wire T138;
  reg [2:0] R139;
  wire[2:0] T140;
  wire T141;
  wire[3:0] T142;
  wire[3:0] idxPagesOH_1;
  wire[3:0] T143;
  wire[1:0] T144;
  wire[1:0] T145;
  wire T146;
  wire[3:0] T147;
  wire[3:0] idxPagesOH_2;
  wire[3:0] T148;
  wire[1:0] T149;
  wire T150;
  wire[3:0] T151;
  wire[3:0] idxPagesOH_3;
  wire[3:0] T152;
  wire[1:0] T153;
  wire[3:0] T154;
  wire[1:0] T155;
  wire T156;
  wire[3:0] T157;
  wire[3:0] idxPagesOH_4;
  wire[3:0] T158;
  wire[1:0] T159;
  wire T160;
  wire[3:0] T161;
  wire[3:0] idxPagesOH_5;
  wire[3:0] T162;
  wire[1:0] T163;
  wire[1:0] T164;
  wire T165;
  wire[3:0] T166;
  wire[3:0] idxPagesOH_6;
  wire[3:0] T167;
  wire[1:0] T168;
  wire T169;
  wire[3:0] T170;
  wire[3:0] idxPagesOH_7;
  wire[3:0] T171;
  wire[1:0] T172;
  wire[7:0] T173;
  wire[7:0] T174;
  wire[7:0] T175;
  wire[3:0] T176;
  wire[1:0] T177;
  wire T178;
  wire[12:0] T179;
  wire[12:0] T180;
  reg [12:0] idxs [7:0];
  wire[12:0] T181;
  wire[12:0] T424;
  wire T182;
  wire[12:0] T183;
  wire[1:0] T184;
  wire T185;
  wire[12:0] T186;
  wire T187;
  wire[12:0] T188;
  wire[3:0] T189;
  wire[1:0] T190;
  wire T191;
  wire[12:0] T192;
  wire T193;
  wire[12:0] T194;
  wire[1:0] T195;
  wire T196;
  wire[12:0] T197;
  wire T198;
  wire[12:0] T199;
  reg [7:0] idxValid;
  wire[7:0] T425;
  wire[7:0] T200;
  wire[7:0] T201;
  wire[7:0] T202;
  wire[7:0] T203;
  wire[7:0] T204;
  wire[7:0] T205;
  wire[7:0] T206;
  wire[3:0] T207;
  wire[1:0] T208;
  wire T209;
  wire[3:0] T210;
  wire[3:0] T211;
  wire[3:0] tgtPagesOH_0;
  wire[3:0] T212;
  wire[1:0] T213;
  reg [1:0] tgtPages [7:0];
  wire[1:0] T214;
  wire[1:0] T426;
  wire T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[3:0] T215;
  wire[1:0] T430;
  wire T431;
  wire T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] tgtPagesOH_1;
  wire[3:0] T219;
  wire[1:0] T220;
  wire[1:0] T221;
  wire T222;
  wire[3:0] T223;
  wire[3:0] T224;
  wire[3:0] tgtPagesOH_2;
  wire[3:0] T225;
  wire[1:0] T226;
  wire T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[3:0] tgtPagesOH_3;
  wire[3:0] T230;
  wire[1:0] T231;
  wire[3:0] T232;
  wire[1:0] T233;
  wire T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] tgtPagesOH_4;
  wire[3:0] T237;
  wire[1:0] T238;
  wire T239;
  wire[3:0] T240;
  wire[3:0] T241;
  wire[3:0] tgtPagesOH_5;
  wire[3:0] T242;
  wire[1:0] T243;
  wire[1:0] T244;
  wire T245;
  wire[3:0] T246;
  wire[3:0] T247;
  wire[3:0] tgtPagesOH_6;
  wire[3:0] T248;
  wire[1:0] T249;
  wire T250;
  wire[3:0] T251;
  wire[3:0] T252;
  wire[3:0] tgtPagesOH_7;
  wire[3:0] T253;
  wire[1:0] T254;
  wire[7:0] T255;
  wire[7:0] T256;
  wire[7:0] T257;
  wire[7:0] T258;
  wire[7:0] T259;
  wire[7:0] T432;
  wire T260;
  wire T261;
  wire[7:0] T262;
  wire[7:0] T263;
  wire[3:0] T433;
  wire[1:0] T434;
  wire T435;
  wire T436;
  wire[42:0] T264;
  wire[42:0] T265;
  wire[42:0] T266;
  wire[12:0] T267;
  wire[12:0] T268;
  wire[12:0] T269;
  reg [12:0] tgts [7:0];
  wire[12:0] T270;
  wire[12:0] T437;
  wire T271;
  wire[12:0] T272;
  wire[12:0] T273;
  wire[12:0] T274;
  wire T275;
  wire[12:0] T276;
  wire[12:0] T277;
  wire[12:0] T278;
  wire T279;
  wire[12:0] T280;
  wire[12:0] T281;
  wire[12:0] T282;
  wire T283;
  wire[12:0] T284;
  wire[12:0] T285;
  wire[12:0] T286;
  wire T287;
  wire[12:0] T288;
  wire[12:0] T289;
  wire[12:0] T290;
  wire T291;
  wire[12:0] T292;
  wire[12:0] T293;
  wire[12:0] T294;
  wire T295;
  wire[12:0] T296;
  wire[12:0] T297;
  wire T298;
  wire[29:0] T299;
  wire[29:0] T300;
  wire[29:0] T301;
  wire T302;
  wire[3:0] T303;
  wire[3:0] T304;
  wire T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire T308;
  wire[3:0] T309;
  wire[3:0] T310;
  wire T311;
  wire[3:0] T312;
  wire[3:0] T313;
  wire T314;
  wire[3:0] T315;
  wire[3:0] T316;
  wire T317;
  wire[3:0] T318;
  wire[3:0] T319;
  wire T320;
  wire[3:0] T321;
  wire[3:0] T322;
  wire T323;
  wire[3:0] T324;
  wire T325;
  wire[29:0] T326;
  wire[29:0] T327;
  wire[29:0] T328;
  wire T329;
  wire[29:0] T330;
  wire[29:0] T331;
  wire[29:0] T332;
  wire T333;
  wire[29:0] T334;
  wire[29:0] T335;
  wire T336;
  wire[42:0] T337;
  reg [42:0] R338;
  wire[42:0] T339;
  wire T340;
  wire T341;
  wire[1:0] T342;
  wire T343;
  wire T344;
  reg  R345;
  wire T438;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  reg [1:0] R352;
  wire[1:0] T439;
  wire[1:0] T353;
  wire[1:0] T354;
  wire[1:0] T355;
  wire[1:0] T356;
  wire T357;
  wire T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  reg [42:0] R365;
  wire[42:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[7:0] T372;
  reg [7:0] useRAS;
  wire[7:0] T373;
  wire[7:0] T374;
  wire[7:0] T375;
  wire[7:0] T376;
  wire[7:0] T377;
  wire[7:0] T378;
  wire[7:0] T440;
  wire T379;
  wire T380;
  reg  R381;
  wire T382;
  wire[7:0] T383;
  wire[7:0] T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire[7:0] T392;
  reg [7:0] isJump;
  wire[7:0] T393;
  wire[7:0] T394;
  wire[7:0] T395;
  wire[7:0] T396;
  wire[7:0] T397;
  wire[7:0] T398;
  wire[7:0] T441;
  wire T399;
  wire T400;
  wire[7:0] T401;
  wire[7:0] T402;
  wire T403;
  wire T404;
  wire T405;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R4 = {2{$random}};
    R8 = {1{$random}};
    updateHit = {1{$random}};
    R15 = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      T18[initvar] = {1{$random}};
    R25 = {1{$random}};
    R31 = {1{$random}};
    R35 = {1{$random}};
    R38 = {1{$random}};
    R42 = {1{$random}};
    pageValid = {1{$random}};
    R62 = {1{$random}};
    R72 = {2{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    R133 = {1{$random}};
    R139 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R338 = {2{$random}};
    R345 = {1{$random}};
    R352 = {1{$random}};
    R365 = {2{$random}};
    useRAS = {1{$random}};
    R381 = {1{$random}};
    isJump = {1{$random}};
  end
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req == R4;
  assign T5 = io_update_valid ? io_update_bits_target : R4;
  assign T6 = T7 ^ 1'h1;
  assign T7 = T11 & updateTarget;
  assign updateTarget = updateValid & R8;
  assign T9 = io_update_valid ? io_update_bits_incorrectTarget : R8;
  assign updateValid = R8 | updateHit;
  assign T10 = io_update_valid ? io_update_bits_prediction_valid : updateHit;
  assign T11 = R15 & T12;
  assign T12 = T13 ^ 1'h1;
  assign T13 = updateValid & T14;
  assign T14 = updateTarget ^ 1'h1;
  assign T406 = reset ? 1'h0 : io_update_valid;
  assign io_resp_bits_bht_value = T16;
  assign T16 = T17;
  assign T17 = T18[T40];
  assign T20 = {R31, T21};
  assign T21 = T28 | T22;
  assign T22 = T23 & R31;
  assign T23 = T27 | T24;
  assign T24 = R25[1'h0:1'h0];
  assign T26 = io_update_valid ? io_update_bits_prediction_bits_bht_value : R25;
  assign T27 = R25[1'h1:1'h1];
  assign T28 = T30 & T29;
  assign T29 = R25[1'h0:1'h0];
  assign T30 = R25[1'h1:1'h1];
  assign T32 = io_update_valid ? io_update_bits_taken : R31;
  assign T33 = T37 & T34;
  assign T34 = R35 ^ 1'h1;
  assign T36 = io_update_valid ? io_update_bits_isJump : R35;
  assign T37 = R15 & updateHit;
  assign T39 = io_update_valid ? io_update_bits_prediction_bits_bht_index : R38;
  assign T40 = T41;
  assign T41 = T46 ^ R42;
  assign T43 = T33 ? T44 : R42;
  assign T44 = {R31, T45};
  assign T45 = R42[2'h3:1'h1];
  assign T46 = io_req[3'h5:2'h2];
  assign io_resp_bits_bht_index = T40;
  assign io_resp_bits_entry = T407;
  assign T407 = {T436, T408};
  assign T408 = {T435, T409};
  assign T409 = T410[1'h1:1'h1];
  assign T410 = T434 | T411;
  assign T411 = T412[1'h1:1'h0];
  assign T412 = T433 | T413;
  assign T413 = hits[2'h3:1'h0];
  assign hits = T173 & T48;
  assign T48 = T49;
  assign T49 = {T154, T50};
  assign T50 = {T145, T51};
  assign T51 = {T141, T52};
  assign T52 = T53 != 4'h0;
  assign T53 = idxPagesOH_0 & pageHit;
  assign pageHit = T116 & pageValid;
  assign T414 = reset ? 4'h0 : T54;
  assign T54 = io_invalidate ? 4'h0 : T55;
  assign T55 = T115 ? T56 : pageValid;
  assign T56 = pageValid | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 4'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T57;
  assign T57 = T59 | T415;
  assign T415 = {3'h0, T58};
  assign T58 = idxPageUpdateOH[2'h3:2'h3];
  assign T59 = T60 << 1'h1;
  assign T60 = idxPageUpdateOH[2'h2:1'h0];
  assign idxPageUpdateOH = useUpdatePageHit ? updatePageHit : idxPageRepl;
  assign idxPageRepl = T61;
  assign T61 = 1'h1 << R62;
  assign T416 = reset ? 2'h0 : T63;
  assign T63 = T65 ? T64 : R62;
  assign T64 = R62 + 2'h1;
  assign T65 = R15 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doIdxPageRepl = updateTarget & T66;
  assign T66 = useUpdatePageHit ^ 1'h1;
  assign updatePageHit = T67 & pageValid;
  assign T67 = T68;
  assign T68 = {T103, T69};
  assign T69 = {T101, T70};
  assign T70 = T74 == T71;
  assign T71 = R72 >> 4'hd;
  assign T73 = io_update_valid ? io_update_bits_pc : R72;
  assign T74 = pages[2'h0];
  assign T76 = T79 ? T78 : T77;
  assign T77 = R72 >> 4'hd;
  assign T78 = io_req >> 4'hd;
  assign T79 = T80 != 4'h0;
  assign T80 = idxPageUpdateOH & 4'h5;
  assign T81 = T11 & T82;
  assign T82 = T84 & T83;
  assign T83 = pageReplEn[2'h3:2'h3];
  assign T84 = T79 ? doTgtPageRepl : doIdxPageRepl;
  assign T86 = T11 & T87;
  assign T87 = T84 & T88;
  assign T88 = pageReplEn[1'h1:1'h1];
  assign T90 = T79 ? T92 : T91;
  assign T91 = io_req >> 4'hd;
  assign T92 = R72 >> 4'hd;
  assign T93 = T11 & T94;
  assign T94 = T96 & T95;
  assign T95 = pageReplEn[2'h2:2'h2];
  assign T96 = T79 ? doIdxPageRepl : doTgtPageRepl;
  assign T98 = T11 & T99;
  assign T99 = T96 & T100;
  assign T100 = pageReplEn[1'h0:1'h0];
  assign T101 = T102 == T71;
  assign T102 = pages[2'h1];
  assign T103 = {T106, T104};
  assign T104 = T105 == T71;
  assign T105 = pages[2'h2];
  assign T106 = T107 == T71;
  assign T107 = pages[2'h3];
  assign useUpdatePageHit = updatePageHit != 4'h0;
  assign samePage = T109 == T108;
  assign T108 = io_req >> 4'hd;
  assign T109 = R72 >> 4'hd;
  assign doTgtPageRepl = T113 & T110;
  assign T110 = usePageHit ^ 1'h1;
  assign usePageHit = T111 != 4'h0;
  assign T111 = pageHit & T112;
  assign T112 = ~ idxPageReplEn;
  assign T113 = updateTarget & T114;
  assign T114 = samePage ^ 1'h1;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 4'h0;
  assign T115 = T11 & doPageRepl;
  assign T116 = T117;
  assign T117 = {T124, T118};
  assign T118 = {T122, T119};
  assign T119 = T121 == T120;
  assign T120 = io_req >> 4'hd;
  assign T121 = pages[2'h0];
  assign T122 = T123 == T120;
  assign T123 = pages[2'h1];
  assign T124 = {T127, T125};
  assign T125 = T126 == T120;
  assign T126 = pages[2'h2];
  assign T127 = T128 == T120;
  assign T128 = pages[2'h3];
  assign idxPagesOH_0 = T129[2'h3:1'h0];
  assign T129 = 1'h1 << T130;
  assign T130 = idxPages[3'h0];
  assign T417 = {T422, T418};
  assign T418 = T419[1'h1:1'h1];
  assign T419 = T421 | T420;
  assign T420 = idxPageUpdateOH[1'h1:1'h0];
  assign T421 = idxPageUpdateOH[2'h3:2'h2];
  assign T422 = T421 != 2'h0;
  assign T132 = updateHit ? R139 : R133;
  assign T423 = reset ? 3'h0 : T134;
  assign T134 = T136 ? T135 : R133;
  assign T135 = R133 + 3'h1;
  assign T136 = T11 & T137;
  assign T137 = T138 & updateValid;
  assign T138 = updateHit ^ 1'h1;
  assign T140 = io_update_valid ? io_update_bits_prediction_bits_entry : R139;
  assign T141 = T142 != 4'h0;
  assign T142 = idxPagesOH_1 & pageHit;
  assign idxPagesOH_1 = T143[2'h3:1'h0];
  assign T143 = 1'h1 << T144;
  assign T144 = idxPages[3'h1];
  assign T145 = {T150, T146};
  assign T146 = T147 != 4'h0;
  assign T147 = idxPagesOH_2 & pageHit;
  assign idxPagesOH_2 = T148[2'h3:1'h0];
  assign T148 = 1'h1 << T149;
  assign T149 = idxPages[3'h2];
  assign T150 = T151 != 4'h0;
  assign T151 = idxPagesOH_3 & pageHit;
  assign idxPagesOH_3 = T152[2'h3:1'h0];
  assign T152 = 1'h1 << T153;
  assign T153 = idxPages[3'h3];
  assign T154 = {T164, T155};
  assign T155 = {T160, T156};
  assign T156 = T157 != 4'h0;
  assign T157 = idxPagesOH_4 & pageHit;
  assign idxPagesOH_4 = T158[2'h3:1'h0];
  assign T158 = 1'h1 << T159;
  assign T159 = idxPages[3'h4];
  assign T160 = T161 != 4'h0;
  assign T161 = idxPagesOH_5 & pageHit;
  assign idxPagesOH_5 = T162[2'h3:1'h0];
  assign T162 = 1'h1 << T163;
  assign T163 = idxPages[3'h5];
  assign T164 = {T169, T165};
  assign T165 = T166 != 4'h0;
  assign T166 = idxPagesOH_6 & pageHit;
  assign idxPagesOH_6 = T167[2'h3:1'h0];
  assign T167 = 1'h1 << T168;
  assign T168 = idxPages[3'h6];
  assign T169 = T170 != 4'h0;
  assign T170 = idxPagesOH_7 & pageHit;
  assign idxPagesOH_7 = T171[2'h3:1'h0];
  assign T171 = 1'h1 << T172;
  assign T172 = idxPages[3'h7];
  assign T173 = idxValid & T174;
  assign T174 = T175;
  assign T175 = {T189, T176};
  assign T176 = {T184, T177};
  assign T177 = {T182, T178};
  assign T178 = T180 == T179;
  assign T179 = io_req[4'hc:1'h0];
  assign T180 = idxs[3'h0];
  assign T424 = R72[4'hc:1'h0];
  assign T182 = T183 == T179;
  assign T183 = idxs[3'h1];
  assign T184 = {T187, T185};
  assign T185 = T186 == T179;
  assign T186 = idxs[3'h2];
  assign T187 = T188 == T179;
  assign T188 = idxs[3'h3];
  assign T189 = {T195, T190};
  assign T190 = {T193, T191};
  assign T191 = T192 == T179;
  assign T192 = idxs[3'h4];
  assign T193 = T194 == T179;
  assign T194 = idxs[3'h5];
  assign T195 = {T198, T196};
  assign T196 = T197 == T179;
  assign T197 = idxs[3'h6];
  assign T198 = T199 == T179;
  assign T199 = idxs[3'h7];
  assign T425 = reset ? 8'h0 : T200;
  assign T200 = io_invalidate ? 8'h0 : T201;
  assign T201 = T11 ? T255 : T202;
  assign T202 = T11 ? T203 : idxValid;
  assign T203 = idxValid & T204;
  assign T204 = ~ T205;
  assign T205 = T206;
  assign T206 = {T232, T207};
  assign T207 = {T221, T208};
  assign T208 = {T216, T209};
  assign T209 = T210 != 4'h0;
  assign T210 = pageReplEn & T211;
  assign T211 = idxPagesOH_0 | tgtPagesOH_0;
  assign tgtPagesOH_0 = T212[2'h3:1'h0];
  assign T212 = 1'h1 << T213;
  assign T213 = tgtPages[3'h0];
  assign T426 = {T431, T427};
  assign T427 = T428[1'h1:1'h1];
  assign T428 = T430 | T429;
  assign T429 = T215[1'h1:1'h0];
  assign T215 = usePageHit ? pageHit : tgtPageRepl;
  assign T430 = T215[2'h3:2'h2];
  assign T431 = T430 != 2'h0;
  assign T216 = T217 != 4'h0;
  assign T217 = pageReplEn & T218;
  assign T218 = idxPagesOH_1 | tgtPagesOH_1;
  assign tgtPagesOH_1 = T219[2'h3:1'h0];
  assign T219 = 1'h1 << T220;
  assign T220 = tgtPages[3'h1];
  assign T221 = {T227, T222};
  assign T222 = T223 != 4'h0;
  assign T223 = pageReplEn & T224;
  assign T224 = idxPagesOH_2 | tgtPagesOH_2;
  assign tgtPagesOH_2 = T225[2'h3:1'h0];
  assign T225 = 1'h1 << T226;
  assign T226 = tgtPages[3'h2];
  assign T227 = T228 != 4'h0;
  assign T228 = pageReplEn & T229;
  assign T229 = idxPagesOH_3 | tgtPagesOH_3;
  assign tgtPagesOH_3 = T230[2'h3:1'h0];
  assign T230 = 1'h1 << T231;
  assign T231 = tgtPages[3'h3];
  assign T232 = {T244, T233};
  assign T233 = {T239, T234};
  assign T234 = T235 != 4'h0;
  assign T235 = pageReplEn & T236;
  assign T236 = idxPagesOH_4 | tgtPagesOH_4;
  assign tgtPagesOH_4 = T237[2'h3:1'h0];
  assign T237 = 1'h1 << T238;
  assign T238 = tgtPages[3'h4];
  assign T239 = T240 != 4'h0;
  assign T240 = pageReplEn & T241;
  assign T241 = idxPagesOH_5 | tgtPagesOH_5;
  assign tgtPagesOH_5 = T242[2'h3:1'h0];
  assign T242 = 1'h1 << T243;
  assign T243 = tgtPages[3'h5];
  assign T244 = {T250, T245};
  assign T245 = T246 != 4'h0;
  assign T246 = pageReplEn & T247;
  assign T247 = idxPagesOH_6 | tgtPagesOH_6;
  assign tgtPagesOH_6 = T248[2'h3:1'h0];
  assign T248 = 1'h1 << T249;
  assign T249 = tgtPages[3'h6];
  assign T250 = T251 != 4'h0;
  assign T251 = pageReplEn & T252;
  assign T252 = idxPagesOH_7 | tgtPagesOH_7;
  assign tgtPagesOH_7 = T253[2'h3:1'h0];
  assign T253 = 1'h1 << T254;
  assign T254 = tgtPages[3'h7];
  assign T255 = T262 | T256;
  assign T256 = T432 & T257;
  assign T257 = T259 | T258;
  assign T258 = idxValid ^ idxValid;
  assign T259 = 1'h1 << T132;
  assign T432 = T260 ? 8'hff : 8'h0;
  assign T260 = T261;
  assign T261 = updateValid;
  assign T262 = T202 & T263;
  assign T263 = ~ T257;
  assign T433 = hits[3'h7:3'h4];
  assign T434 = T412[2'h3:2'h2];
  assign T435 = T434 != 2'h0;
  assign T436 = T433 != 4'h0;
  assign io_resp_bits_target = T264;
  assign T264 = T387 ? io_update_bits_returnAddr : T265;
  assign T265 = T370 ? T337 : T266;
  assign T266 = {T299, T267};
  assign T267 = T272 | T268;
  assign T268 = T271 ? T269 : 13'h0;
  assign T269 = tgts[3'h7];
  assign T437 = io_req[4'hc:1'h0];
  assign T271 = hits[3'h7:3'h7];
  assign T272 = T276 | T273;
  assign T273 = T275 ? T274 : 13'h0;
  assign T274 = tgts[3'h6];
  assign T275 = hits[3'h6:3'h6];
  assign T276 = T280 | T277;
  assign T277 = T279 ? T278 : 13'h0;
  assign T278 = tgts[3'h5];
  assign T279 = hits[3'h5:3'h5];
  assign T280 = T284 | T281;
  assign T281 = T283 ? T282 : 13'h0;
  assign T282 = tgts[3'h4];
  assign T283 = hits[3'h4:3'h4];
  assign T284 = T288 | T285;
  assign T285 = T287 ? T286 : 13'h0;
  assign T286 = tgts[3'h3];
  assign T287 = hits[2'h3:2'h3];
  assign T288 = T292 | T289;
  assign T289 = T291 ? T290 : 13'h0;
  assign T290 = tgts[3'h2];
  assign T291 = hits[2'h2:2'h2];
  assign T292 = T296 | T293;
  assign T293 = T295 ? T294 : 13'h0;
  assign T294 = tgts[3'h1];
  assign T295 = hits[1'h1:1'h1];
  assign T296 = T298 ? T297 : 13'h0;
  assign T297 = tgts[3'h0];
  assign T298 = hits[1'h0:1'h0];
  assign T299 = T326 | T300;
  assign T300 = T302 ? T301 : 30'h0;
  assign T301 = pages[2'h3];
  assign T302 = T303[2'h3:2'h3];
  assign T303 = T306 | T304;
  assign T304 = T305 ? tgtPagesOH_7 : 4'h0;
  assign T305 = hits[3'h7:3'h7];
  assign T306 = T309 | T307;
  assign T307 = T308 ? tgtPagesOH_6 : 4'h0;
  assign T308 = hits[3'h6:3'h6];
  assign T309 = T312 | T310;
  assign T310 = T311 ? tgtPagesOH_5 : 4'h0;
  assign T311 = hits[3'h5:3'h5];
  assign T312 = T315 | T313;
  assign T313 = T314 ? tgtPagesOH_4 : 4'h0;
  assign T314 = hits[3'h4:3'h4];
  assign T315 = T318 | T316;
  assign T316 = T317 ? tgtPagesOH_3 : 4'h0;
  assign T317 = hits[2'h3:2'h3];
  assign T318 = T321 | T319;
  assign T319 = T320 ? tgtPagesOH_2 : 4'h0;
  assign T320 = hits[2'h2:2'h2];
  assign T321 = T324 | T322;
  assign T322 = T323 ? tgtPagesOH_1 : 4'h0;
  assign T323 = hits[1'h1:1'h1];
  assign T324 = T325 ? tgtPagesOH_0 : 4'h0;
  assign T325 = hits[1'h0:1'h0];
  assign T326 = T330 | T327;
  assign T327 = T329 ? T328 : 30'h0;
  assign T328 = pages[2'h2];
  assign T329 = T303[2'h2:2'h2];
  assign T330 = T334 | T331;
  assign T331 = T333 ? T332 : 30'h0;
  assign T332 = pages[2'h1];
  assign T333 = T303[1'h1:1'h1];
  assign T334 = T336 ? T335 : 30'h0;
  assign T335 = pages[2'h0];
  assign T336 = T303[1'h0:1'h0];
  assign T337 = T369 ? R365 : R338;
  assign T339 = T340 ? io_update_bits_returnAddr : R338;
  assign T340 = T364 & T341;
  assign T341 = T342[1'h0:1'h0];
  assign T342 = 1'h1 << T343;
  assign T343 = T344;
  assign T344 = R345 + 1'h1;
  assign T438 = reset ? 1'h0 : T346;
  assign T346 = T349 ? T348 : T347;
  assign T347 = T364 ? T344 : R345;
  assign T348 = R345 - 1'h1;
  assign T349 = T360 & T350;
  assign T350 = T351 ^ 1'h1;
  assign T351 = R352 == 2'h0;
  assign T439 = reset ? 2'h0 : T353;
  assign T353 = io_invalidate ? 2'h0 : T354;
  assign T354 = T349 ? T359 : T355;
  assign T355 = T357 ? T356 : R352;
  assign T356 = R352 + 2'h1;
  assign T357 = T364 & T358;
  assign T358 = R352 < 2'h2;
  assign T359 = R352 - 2'h1;
  assign T360 = io_update_valid & T361;
  assign T361 = T363 & T362;
  assign T362 = io_update_bits_isReturn & io_update_bits_prediction_valid;
  assign T363 = io_update_bits_isCall ^ 1'h1;
  assign T364 = io_update_valid & io_update_bits_isCall;
  assign T366 = T367 ? io_update_bits_returnAddr : R365;
  assign T367 = T364 & T368;
  assign T368 = T342[1'h1:1'h1];
  assign T369 = R345;
  assign T370 = T385 & T371;
  assign T371 = T372 != 8'h0;
  assign T372 = hits & useRAS;
  assign T373 = T7 ? T374 : useRAS;
  assign T374 = T383 | T375;
  assign T375 = T440 & T376;
  assign T376 = T378 | T377;
  assign T377 = useRAS ^ useRAS;
  assign T378 = 1'h1 << T132;
  assign T440 = T379 ? 8'hff : 8'h0;
  assign T379 = T380;
  assign T380 = R381;
  assign T382 = io_update_valid ? io_update_bits_isReturn : R381;
  assign T383 = useRAS & T384;
  assign T384 = ~ T376;
  assign T385 = T386 ^ 1'h1;
  assign T386 = R352 == 2'h0;
  assign T387 = T364 & T371;
  assign io_resp_bits_taken = T388;
  assign T388 = T389 ? 1'h0 : io_resp_valid;
  assign T389 = T403 & T390;
  assign T390 = T391 ^ 1'h1;
  assign T391 = T392 != 8'h0;
  assign T392 = hits & isJump;
  assign T393 = T7 ? T394 : isJump;
  assign T394 = T401 | T395;
  assign T395 = T441 & T396;
  assign T396 = T398 | T397;
  assign T397 = isJump ^ isJump;
  assign T398 = 1'h1 << T132;
  assign T441 = T399 ? 8'hff : 8'h0;
  assign T399 = T400;
  assign T400 = R35;
  assign T401 = isJump & T402;
  assign T402 = ~ T396;
  assign T403 = T404 ^ 1'h1;
  assign T404 = T16[1'h0:1'h0];
  assign io_resp_valid = T405;
  assign T405 = hits != 8'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
`endif
    if(io_update_valid) begin
      R4 <= io_update_bits_target;
    end
    if(io_update_valid) begin
      R8 <= io_update_bits_incorrectTarget;
    end
    if(io_update_valid) begin
      updateHit <= io_update_bits_prediction_valid;
    end
    if(reset) begin
      R15 <= 1'h0;
    end else begin
      R15 <= io_update_valid;
    end
    if (T33)
      T18[R38] <= T20;
    if(io_update_valid) begin
      R25 <= io_update_bits_prediction_bits_bht_value;
    end
    if(io_update_valid) begin
      R31 <= io_update_bits_taken;
    end
    if(io_update_valid) begin
      R35 <= io_update_bits_isJump;
    end
    if(io_update_valid) begin
      R38 <= io_update_bits_prediction_bits_bht_index;
    end
    if(T33) begin
      R42 <= T44;
    end
    if(reset) begin
      pageValid <= 4'h0;
    end else if(io_invalidate) begin
      pageValid <= 4'h0;
    end else if(T115) begin
      pageValid <= T56;
    end
    if(reset) begin
      R62 <= 2'h0;
    end else if(T65) begin
      R62 <= T64;
    end
    if(io_update_valid) begin
      R72 <= io_update_bits_pc;
    end
    if (T81)
      pages[2'h3] <= T76;
    if (T86)
      pages[2'h1] <= T76;
    if (T93)
      pages[2'h2] <= T90;
    if (T98)
      pages[2'h0] <= T90;
    if (T7)
      idxPages[T132] <= T417;
    if(reset) begin
      R133 <= 3'h0;
    end else if(T136) begin
      R133 <= T135;
    end
    if(io_update_valid) begin
      R139 <= io_update_bits_prediction_bits_entry;
    end
    if (T7)
      idxs[T132] <= T424;
    if(reset) begin
      idxValid <= 8'h0;
    end else if(io_invalidate) begin
      idxValid <= 8'h0;
    end else if(T11) begin
      idxValid <= T255;
    end else if(T11) begin
      idxValid <= T203;
    end
    if (T7)
      tgtPages[T132] <= T426;
    if (T7)
      tgts[T132] <= T437;
    if(T340) begin
      R338 <= io_update_bits_returnAddr;
    end
    if(reset) begin
      R345 <= 1'h0;
    end else if(T349) begin
      R345 <= T348;
    end else if(T364) begin
      R345 <= T344;
    end
    if(reset) begin
      R352 <= 2'h0;
    end else if(io_invalidate) begin
      R352 <= 2'h0;
    end else if(T349) begin
      R352 <= T359;
    end else if(T357) begin
      R352 <= T356;
    end
    if(T367) begin
      R365 <= io_update_bits_returnAddr;
    end
    if(T7) begin
      useRAS <= T374;
    end
    if(io_update_valid) begin
      R381 <= io_update_bits_isReturn;
    end
    if(T7) begin
      isJump <= T394;
    end
  end
endmodule

module FlowThroughSerializer_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [1:0] io_in_bits_payload_client_xact_id,
    input [2:0] io_in_bits_payload_master_xact_id,
    input [3:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T36;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T37;
  wire T4;
  wire T5;
  reg  active;
  wire T38;
  wire T6;
  wire T7;
  wire[1:0] T8;
  wire T9;
  wire[3:0] T10;
  reg [3:0] rbits_payload_g_type;
  wire[3:0] T39;
  wire[3:0] T11;
  wire[2:0] T12;
  reg [2:0] rbits_payload_master_xact_id;
  wire[2:0] T40;
  wire[2:0] T13;
  wire[1:0] T14;
  reg [1:0] rbits_payload_client_xact_id;
  wire[1:0] T41;
  wire[1:0] T15;
  wire[511:0] T16;
  wire[511:0] T17;
  reg [511:0] rbits_payload_data;
  wire[511:0] T42;
  wire[511:0] T18;
  wire[511:0] T43;
  wire[127:0] T19;
  wire[127:0] T20;
  wire[127:0] shifter_0;
  wire[127:0] T21;
  wire[127:0] shifter_1;
  wire[127:0] T22;
  wire T23;
  wire[1:0] T24;
  wire[127:0] T25;
  wire[127:0] shifter_2;
  wire[127:0] T26;
  wire[127:0] shifter_3;
  wire[127:0] T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  reg [1:0] rbits_header_dst;
  wire[1:0] T44;
  wire[1:0] T31;
  wire[1:0] T32;
  reg [1:0] rbits_header_src;
  wire[1:0] T45;
  wire[1:0] T33;
  wire T34;
  wire T35;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cnt = {1{$random}};
    active = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T9 & wrap;
  assign wrap = cnt == 2'h3;
  assign T36 = reset ? 2'h0 : T1;
  assign T1 = T0 ? 2'h0 : T2;
  assign T2 = T9 ? T8 : T3;
  assign T3 = T4 ? T37 : cnt;
  assign T37 = {1'h0, io_out_ready};
  assign T4 = T5 & io_in_valid;
  assign T5 = active ^ 1'h1;
  assign T38 = reset ? 1'h0 : T6;
  assign T6 = T0 ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : active;
  assign T8 = cnt + 2'h1;
  assign T9 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T10;
  assign T10 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T39 = reset ? io_in_bits_payload_g_type : T11;
  assign T11 = T4 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_master_xact_id = T12;
  assign T12 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T40 = reset ? io_in_bits_payload_master_xact_id : T13;
  assign T13 = T4 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T14;
  assign T14 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T41 = reset ? io_in_bits_payload_client_xact_id : T15;
  assign T15 = T4 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T16;
  assign T16 = active ? T43 : T17;
  assign T17 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T42 = reset ? io_in_bits_payload_data : T18;
  assign T18 = T4 ? io_in_bits_payload_data : rbits_payload_data;
  assign T43 = {384'h0, T19};
  assign T19 = T29 ? T25 : T20;
  assign T20 = T23 ? shifter_1 : shifter_0;
  assign shifter_0 = T21;
  assign T21 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T22;
  assign T22 = rbits_payload_data[8'hff:8'h80];
  assign T23 = T24[1'h0:1'h0];
  assign T24 = cnt;
  assign T25 = T28 ? shifter_3 : shifter_2;
  assign shifter_2 = T26;
  assign T26 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T27;
  assign T27 = rbits_payload_data[9'h1ff:9'h180];
  assign T28 = T24[1'h0:1'h0];
  assign T29 = T24[1'h1:1'h1];
  assign io_out_bits_header_dst = T30;
  assign T30 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T44 = reset ? io_in_bits_header_dst : T31;
  assign T31 = T4 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T32;
  assign T32 = active ? rbits_header_src : io_in_bits_header_src;
  assign T45 = reset ? io_in_bits_header_src : T33;
  assign T33 = T4 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T34;
  assign T34 = active | io_in_valid;
  assign io_in_ready = T35;
  assign T35 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      cnt <= 2'h0;
    end else if(T0) begin
      cnt <= 2'h0;
    end else if(T9) begin
      cnt <= T8;
    end else if(T4) begin
      cnt <= T37;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T0) begin
      active <= 1'h0;
    end else if(T4) begin
      active <= 1'h1;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T4) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T4) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T4) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T4) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T4) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T4) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output io_count
);

  wire T13;
  wire[1:0] T0;
  reg  full;
  wire T14;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[2:0] T3;
  wire[6:0] T4;
  reg [6:0] ram [0:0];
  wire[6:0] T5;
  wire[6:0] T6;
  wire[6:0] T7;
  wire[4:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire empty;
  wire T12;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T13;
  assign T13 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T14 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_master_xact_id = T3;
  assign T3 = T4[2'h2:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {io_enq_bits_header_src, T8};
  assign T8 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign io_deq_bits_header_dst = T9;
  assign T9 = T4[3'h4:2'h3];
  assign io_deq_bits_header_src = T10;
  assign T10 = T4[3'h6:3'h5];
  assign io_deq_valid = T11;
  assign T11 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [12:0] io_req_bits_idx,
    input [18:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[31:0] io_resp_bits_data,
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id
);

  wire T128;
  wire T129;
  wire[3:0] T0;
  wire[2:0] T1;
  wire[5:0] T2;
  wire[2:0] T3;
  wire[511:0] T4;
  wire[1:0] T5;
  wire[25:0] T6;
  wire[25:0] T7;
  reg [31:0] s2_addr;
  wire[31:0] T8;
  wire[31:0] s1_addr;
  wire[31:0] T9;
  reg [12:0] s1_pgoff;
  wire[12:0] T10;
  wire T11;
  wire rdy;
  wire T12;
  wire T13;
  wire s2_miss;
  wire T14;
  wire s2_any_tag_hit;
  wire T15;
  wire T16;
  wire s2_disparity_0;
  wire T17;
  reg  R18;
  wire T19;
  wire T20;
  wire T21;
  wire stall;
  wire T22;
  reg  s1_valid;
  wire T117;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  reg  R28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[6:0] T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[5:0] T37;
  wire T38;
  reg [63:0] vb_array;
  wire[63:0] T118;
  wire[127:0] T119;
  wire[127:0] T39;
  wire[127:0] T40;
  wire[127:0] T41;
  wire[127:0] T120;
  wire[127:0] T42;
  wire[127:0] T43;
  wire[127:0] T44;
  wire[6:0] T45;
  wire[5:0] s2_idx;
  wire[127:0] T121;
  wire T46;
  wire[127:0] T47;
  wire[127:0] T48;
  wire[127:0] T122;
  wire T49;
  wire T50;
  reg  invalidated;
  wire T51;
  wire T52;
  wire T53;
  reg [1:0] state;
  wire[1:0] T123;
  wire[1:0] T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[127:0] T66;
  wire[127:0] T67;
  wire[127:0] T68;
  wire[6:0] T69;
  wire[127:0] T124;
  wire T70;
  wire[127:0] T71;
  wire[127:0] T72;
  wire[127:0] T125;
  wire T73;
  wire s2_tag_hit_0;
  wire T74;
  reg  R75;
  wire T76;
  wire s1_tag_match_0;
  wire T77;
  wire[19:0] s1_tag;
  wire[19:0] T78;
  wire[19:0] T79;
  wire[19:0] T80;
  wire T87;
  wire s0_valid;
  wire T88;
  wire T89;
  wire[5:0] T85;
  wire[12:0] s0_pgoff;
  wire T86;
  wire[19:0] T81;
  wire[19:0] T82;
  wire[19:0] T83;
  wire[19:0] s2_tag;
  reg [5:0] tag_raddr;
  wire[5:0] T84;
  reg  s2_valid;
  wire T126;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [127:0] s2_dout_0;
  wire[127:0] T101;
  wire[127:0] T102;
  wire T109;
  wire T110;
  wire[7:0] T108;
  wire[127:0] T104;
  wire[127:0] T127;
  wire[7:0] T105;
  reg [7:0] R106;
  wire[7:0] T107;
  wire T111;
  wire T112;
  wire T113;
  wire[31:0] s2_dout_word_0;
  wire[127:0] T114;
  wire[6:0] T115;
  wire[1:0] T116;
  wire[5:0] s2_offset;
  wire s2_hit;
  wire FlowThroughSerializer_1_io_in_ready;
  wire FlowThroughSerializer_1_io_out_valid;
  wire[1:0] FlowThroughSerializer_1_io_out_bits_header_src;
  wire[511:0] FlowThroughSerializer_1_io_out_bits_payload_data;
  wire[2:0] FlowThroughSerializer_1_io_out_bits_payload_master_xact_id;
  wire[3:0] FlowThroughSerializer_1_io_out_bits_payload_g_type;
  wire[1:0] FlowThroughSerializer_1_io_cnt;
  wire FlowThroughSerializer_1_io_done;
  wire ack_q_io_enq_ready;
  wire ack_q_io_deq_valid;
  wire[1:0] ack_q_io_deq_bits_header_src;
  wire[1:0] ack_q_io_deq_bits_header_dst;
  wire[2:0] ack_q_io_deq_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_addr = {1{$random}};
    s1_pgoff = {1{$random}};
    R18 = {1{$random}};
    s1_valid = {1{$random}};
    R28 = {1{$random}};
    vb_array = {2{$random}};
    invalidated = {1{$random}};
    state = {1{$random}};
    R75 = {1{$random}};
    tag_raddr = {1{$random}};
    s2_valid = {1{$random}};
    s2_dout_0 = {4{$random}};
    R106 = {1{$random}};
  end
`endif

  assign T128 = FlowThroughSerializer_1_io_done & T129;
  assign T129 = FlowThroughSerializer_1_io_out_bits_payload_g_type != 4'h0;
  assign io_mem_finish_bits_payload_master_xact_id = ack_q_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ack_q_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ack_q_io_deq_bits_header_src;
  assign io_mem_finish_valid = ack_q_io_deq_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_1_io_in_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = T0;
  assign T0 = 4'h0;
  assign io_mem_acquire_bits_payload_subword_addr = T1;
  assign T1 = 3'h0;
  assign io_mem_acquire_bits_payload_write_mask = T2;
  assign T2 = 6'h0;
  assign io_mem_acquire_bits_payload_a_type = T3;
  assign T3 = 3'h2;
  assign io_mem_acquire_bits_payload_data = T4;
  assign T4 = 512'h0;
  assign io_mem_acquire_bits_payload_client_xact_id = T5;
  assign T5 = 2'h0;
  assign io_mem_acquire_bits_payload_addr = T6;
  assign T6 = T7;
  assign T7 = s2_addr >> 3'h6;
  assign T8 = T96 ? s1_addr : s2_addr;
  assign s1_addr = T9;
  assign T9 = {io_req_bits_ppn, s1_pgoff};
  assign T10 = T11 ? io_req_bits_idx : s1_pgoff;
  assign T11 = io_req_valid & rdy;
  assign rdy = T12;
  assign T12 = T95 & T13;
  assign T13 = s2_miss ^ 1'h1;
  assign s2_miss = s2_valid & T14;
  assign T14 = s2_any_tag_hit ^ 1'h1;
  assign s2_any_tag_hit = T15;
  assign T15 = s2_tag_hit_0 & T16;
  assign T16 = s2_disparity_0 ^ 1'h1;
  assign s2_disparity_0 = T17;
  assign T17 = R28 & R18;
  assign T19 = T20 ? 1'h0 : R18;
  assign T20 = T22 & T21;
  assign T21 = stall ^ 1'h1;
  assign stall = io_resp_ready ^ 1'h1;
  assign T22 = s1_valid & rdy;
  assign T117 = reset ? 1'h0 : T23;
  assign T23 = T27 | T24;
  assign T24 = T26 & T25;
  assign T25 = io_req_bits_kill ^ 1'h1;
  assign T26 = s1_valid & stall;
  assign T27 = io_req_valid & rdy;
  assign T29 = T20 ? T30 : R28;
  assign T30 = T31;
  assign T31 = T38 & T32;
  assign T32 = T33 - 1'h1;
  assign T33 = 1'h1 << T34;
  assign T34 = T35 + 7'h1;
  assign T35 = T36 - T36;
  assign T36 = {1'h0, T37};
  assign T37 = s1_pgoff[4'hb:3'h6];
  assign T38 = vb_array >> T36;
  assign T118 = T119[6'h3f:1'h0];
  assign T119 = reset ? 128'h0 : T39;
  assign T39 = T73 ? T66 : T40;
  assign T40 = io_invalidate ? 128'h0 : T41;
  assign T41 = T49 ? T42 : T120;
  assign T120 = {64'h0, vb_array};
  assign T42 = T47 | T43;
  assign T43 = T121 & T44;
  assign T44 = 1'h1 << T45;
  assign T45 = {1'h0, s2_idx};
  assign s2_idx = s2_addr[4'hb:3'h6];
  assign T121 = T46 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T46 = 1'h1;
  assign T47 = T122 & T48;
  assign T48 = ~ T44;
  assign T122 = {64'h0, vb_array};
  assign T49 = FlowThroughSerializer_1_io_done & T50;
  assign T50 = invalidated ^ 1'h1;
  assign T51 = T53 ? 1'h0 : T52;
  assign T52 = io_invalidate ? 1'h1 : invalidated;
  assign T53 = 2'h0 == state;
  assign T123 = reset ? 2'h0 : T54;
  assign T54 = T64 ? 2'h0 : T55;
  assign T55 = T62 ? 2'h3 : T56;
  assign T56 = T59 ? 2'h2 : T57;
  assign T57 = T58 ? 2'h1 : state;
  assign T58 = T53 & s2_miss;
  assign T59 = T61 & T60;
  assign T60 = io_mem_acquire_ready & ack_q_io_enq_ready;
  assign T61 = 2'h1 == state;
  assign T62 = T63 & io_mem_grant_valid;
  assign T63 = 2'h2 == state;
  assign T64 = T65 & FlowThroughSerializer_1_io_done;
  assign T65 = 2'h3 == state;
  assign T66 = T71 | T67;
  assign T67 = T124 & T68;
  assign T68 = 1'h1 << T69;
  assign T69 = {1'h0, s2_idx};
  assign T124 = T70 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T70 = 1'h0;
  assign T71 = T125 & T72;
  assign T72 = ~ T68;
  assign T125 = {64'h0, vb_array};
  assign T73 = s2_valid & s2_disparity_0;
  assign s2_tag_hit_0 = T74;
  assign T74 = R28 & R75;
  assign T76 = T20 ? s1_tag_match_0 : R75;
  assign s1_tag_match_0 = T77;
  assign T77 = T78 == s1_tag;
  assign s1_tag = s1_addr[5'h1f:4'hc];
  assign T78 = T79[5'h13:1'h0];
  assign T79 = T80[5'h13:1'h0];
  assign T87 = T89 & s0_valid;
  assign s0_valid = io_req_valid | T88;
  assign T88 = s1_valid & stall;
  assign T89 = FlowThroughSerializer_1_io_done ^ 1'h1;
  assign T85 = s0_pgoff[4'hb:3'h6];
  assign s0_pgoff = T86 ? s1_pgoff : io_req_bits_idx;
  assign T86 = s1_valid & stall;
  ICache_tag_array tag_array (
    .CLK(clk),
    .RW0A(FlowThroughSerializer_1_io_done ? s2_idx : T85),
    .RW0E(T87 || FlowThroughSerializer_1_io_done),
    .RW0W(FlowThroughSerializer_1_io_done),
    .RW0I(T83),
    .RW0M(T82),
    .RW0O(T80)
  );
  assign T82 = 20'hfffff;
  assign T83 = s2_tag;
  assign s2_tag = s2_addr[5'h1f:4'hc];
  assign T84 = T87 ? T85 : tag_raddr;
  assign T126 = reset ? 1'h0 : T90;
  assign T90 = T92 | T91;
  assign T91 = io_resp_valid & stall;
  assign T92 = T94 & T93;
  assign T93 = io_req_bits_kill ^ 1'h1;
  assign T94 = s1_valid & rdy;
  assign T95 = state == 2'h0;
  assign T96 = T98 & T97;
  assign T97 = stall ^ 1'h1;
  assign T98 = s1_valid & rdy;
  assign io_mem_acquire_valid = T99;
  assign T99 = T100 & ack_q_io_enq_ready;
  assign T100 = state == 2'h1;
  assign io_resp_bits_datablock = s2_dout_0;
  assign T101 = T111 ? T102 : s2_dout_0;
  assign T109 = T110 & s0_valid;
  assign T110 = FlowThroughSerializer_1_io_out_valid ^ 1'h1;
  assign T108 = s0_pgoff[4'hb:3'h4];
  ICache_T103 T103 (
    .CLK(clk),
    .RW0A(FlowThroughSerializer_1_io_out_valid ? T105 : T108),
    .RW0E(T109 || FlowThroughSerializer_1_io_out_valid),
    .RW0W(FlowThroughSerializer_1_io_out_valid),
    .RW0I(T127),
    .RW0O(T102)
  );
  assign T127 = FlowThroughSerializer_1_io_out_bits_payload_data[7'h7f:1'h0];
  assign T105 = {s2_idx, FlowThroughSerializer_1_io_cnt};
  assign T107 = T109 ? T108 : R106;
  assign T111 = T113 & T112;
  assign T112 = stall ^ 1'h1;
  assign T113 = s1_valid & rdy;
  assign io_resp_bits_data = s2_dout_word_0;
  assign s2_dout_word_0 = T114[5'h1f:1'h0];
  assign T114 = s2_dout_0 >> T115;
  assign T115 = T116 << 3'h5;
  assign T116 = s2_offset[2'h3:2'h2];
  assign s2_offset = s2_addr[3'h5:1'h0];
  assign io_resp_valid = s2_hit;
  assign s2_hit = s2_valid & s2_any_tag_hit;
  FlowThroughSerializer_1 FlowThroughSerializer_1(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_1_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( FlowThroughSerializer_1_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_1_io_out_bits_header_src ),
       //.io_out_bits_header_dst(  )
       .io_out_bits_payload_data( FlowThroughSerializer_1_io_out_bits_payload_data ),
       //.io_out_bits_payload_client_xact_id(  )
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_1_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_1_io_out_bits_payload_g_type ),
       .io_cnt( FlowThroughSerializer_1_io_cnt ),
       .io_done( FlowThroughSerializer_1_io_done )
  );
  Queue_11 ack_q(.clk(clk), .reset(reset),
       .io_enq_ready( ack_q_io_enq_ready ),
       .io_enq_valid( T128 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( FlowThroughSerializer_1_io_out_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( FlowThroughSerializer_1_io_out_bits_payload_master_xact_id ),
       .io_deq_ready( io_mem_finish_ready ),
       .io_deq_valid( ack_q_io_deq_valid ),
       .io_deq_bits_header_src( ack_q_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ack_q_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ack_q_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ack_q.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(T96) begin
      s2_addr <= s1_addr;
    end
    if(T11) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(T20) begin
      R18 <= 1'h0;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T23;
    end
    if(T20) begin
      R28 <= T30;
    end
    vb_array <= T118;
    if(T53) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T64) begin
      state <= 2'h0;
    end else if(T62) begin
      state <= 2'h3;
    end else if(T59) begin
      state <= 2'h2;
    end else if(T58) begin
      state <= 2'h1;
    end
    if(T20) begin
      R75 <= s1_tag_match_0;
    end
    if(T87) begin
      tag_raddr <= T85;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= T90;
    end
    if(T111) begin
      s2_dout_0 <= T102;
    end
    if(T109) begin
      R106 <= T108;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input  io_clear_hit,
    input [36:0] io_tag,
    output io_hit,
    output[3:0] io_hits,
    output[3:0] io_valid_bits,
    input  io_write,
    input [36:0] io_write_tag,
    input [1:0] io_write_addr
);

  reg [3:0] vb_array;
  wire[3:0] T31;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T32;
  wire T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire T11;
  wire T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[1:0] T15;
  wire hits_0;
  wire T16;
  wire[36:0] T17;
  reg [36:0] cam_tags [3:0];
  wire[36:0] T18;
  wire T19;
  wire hits_1;
  wire T20;
  wire[36:0] T21;
  wire T22;
  wire[1:0] T23;
  wire hits_2;
  wire T24;
  wire[36:0] T25;
  wire T26;
  wire hits_3;
  wire T27;
  wire[36:0] T28;
  wire T29;
  wire T30;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
`endif

  assign io_valid_bits = vb_array;
  assign T31 = reset ? 4'h0 : T0;
  assign T0 = T11 ? T9 : T1;
  assign T1 = io_clear ? 4'h0 : T2;
  assign T2 = io_write ? T3 : vb_array;
  assign T3 = T7 | T4;
  assign T4 = T32 & T5;
  assign T5 = 1'h1 << io_write_addr;
  assign T32 = T6 ? 4'hf : 4'h0;
  assign T6 = 1'h1;
  assign T7 = vb_array & T8;
  assign T8 = ~ T5;
  assign T9 = vb_array & T10;
  assign T10 = ~ io_hits;
  assign T11 = T12 & io_clear_hit;
  assign T12 = io_clear ^ 1'h1;
  assign io_hits = T13;
  assign T13 = T14;
  assign T14 = {T23, T15};
  assign T15 = {hits_1, hits_0};
  assign hits_0 = T19 & T16;
  assign T16 = T17 == io_tag;
  assign T17 = cam_tags[2'h0];
  assign T19 = vb_array[1'h0:1'h0];
  assign hits_1 = T22 & T20;
  assign T20 = T21 == io_tag;
  assign T21 = cam_tags[2'h1];
  assign T22 = vb_array[1'h1:1'h1];
  assign T23 = {hits_3, hits_2};
  assign hits_2 = T26 & T24;
  assign T24 = T25 == io_tag;
  assign T25 = cam_tags[2'h2];
  assign T26 = vb_array[2'h2:2'h2];
  assign hits_3 = T29 & T27;
  assign T27 = T28 == io_tag;
  assign T28 = cam_tags[2'h3];
  assign T29 = vb_array[2'h3:2'h3];
  assign io_hit = T30;
  assign T30 = io_hits != 4'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 4'h0;
    end else if(T11) begin
      vb_array <= T9;
    end else if(io_clear) begin
      vb_array <= 4'h0;
    end else if(io_write) begin
      vb_array <= T3;
    end
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [30:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    output io_resp_miss,
    output[3:0] io_resp_hit_idx,
    output[18:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[29:0] io_ptw_req_bits,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [18:0] io_ptw_resp_bits_ppn,
    input [5:0] io_ptw_resp_bits_perm,
    input [7:0] io_ptw_status_ip,
    input [7:0] io_ptw_status_im,
    input [6:0] io_ptw_status_zero,
    input  io_ptw_status_er,
    input  io_ptw_status_vm,
    input  io_ptw_status_s64,
    input  io_ptw_status_u64,
    input  io_ptw_status_ef,
    input  io_ptw_status_pei,
    input  io_ptw_status_ei,
    input  io_ptw_status_ps,
    input  io_ptw_status_s,
    input  io_ptw_invalidate,
    input  io_ptw_sret
);

  reg [1:0] r_refill_waddr;
  wire[1:0] T32;
  wire[1:0] repl_waddr;
  wire[1:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire T40;
  reg [3:0] R41;
  wire[3:0] T42;
  wire[3:0] T43;
  wire[3:0] T44;
  wire[3:0] T45;
  wire[6:0] T46;
  wire[1:0] T47;
  wire T48;
  wire[1:0] T149;
  wire T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire T154;
  wire T50;
  wire[3:0] T51;
  wire[3:0] T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire T56;
  wire tlb_hit;
  wire[1:0] T57;
  wire T58;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[1:0] T157;
  wire T158;
  wire[3:0] T59;
  wire T159;
  wire T160;
  wire has_invalid_entry;
  wire T60;
  wire T2;
  wire tlb_miss;
  wire T3;
  wire bad_va;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[36:0] T168;
  reg [37:0] r_refill_tag;
  wire[37:0] T0;
  wire[37:0] lookup_tag;
  wire[37:0] T1;
  wire T169;
  wire T170;
  reg [1:0] state;
  wire[1:0] T148;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[36:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire[29:0] T147;
  wire T9;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] T27;
  reg [3:0] ux_array;
  wire[3:0] T28;
  wire[3:0] T29;
  wire[3:0] T30;
  wire[3:0] T31;
  wire[3:0] T161;
  wire T61;
  wire T62;
  wire[5:0] T63;
  wire[5:0] T162;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire[3:0] T67;
  wire T68;
  wire[3:0] T69;
  reg [3:0] sx_array;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire[3:0] T163;
  wire T74;
  wire T75;
  wire[3:0] T76;
  wire[3:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire[3:0] T83;
  reg [3:0] uw_array;
  wire[3:0] T84;
  wire[3:0] T85;
  wire[3:0] T86;
  wire[3:0] T87;
  wire[3:0] T164;
  wire T88;
  wire T89;
  wire[3:0] T90;
  wire[3:0] T91;
  wire T92;
  wire[3:0] T93;
  reg [3:0] sw_array;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] T97;
  wire[3:0] T165;
  wire T98;
  wire T99;
  wire[3:0] T100;
  wire[3:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire[3:0] T107;
  reg [3:0] ur_array;
  wire[3:0] T108;
  wire[3:0] T109;
  wire[3:0] T110;
  wire[3:0] T111;
  wire[3:0] T166;
  wire T112;
  wire T113;
  wire[3:0] T114;
  wire[3:0] T115;
  wire T116;
  wire[3:0] T117;
  reg [3:0] sr_array;
  wire[3:0] T118;
  wire[3:0] T119;
  wire[3:0] T120;
  wire[3:0] T121;
  wire[3:0] T167;
  wire T122;
  wire T123;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[18:0] T126;
  wire[18:0] T127;
  wire[18:0] T128;
  wire[18:0] T129;
  wire[18:0] T130;
  reg [18:0] tag_ram [3:0];
  wire[18:0] T131;
  wire T132;
  wire[18:0] T133;
  wire[18:0] T134;
  wire[18:0] T135;
  wire T136;
  wire[18:0] T137;
  wire[18:0] T138;
  wire[18:0] T139;
  wire T140;
  wire[18:0] T141;
  wire[18:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire tag_cam_io_hit;
  wire[3:0] tag_cam_io_hits;
  wire[3:0] tag_cam_io_valid_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R41 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    ux_array = {1{$random}};
    sx_array = {1{$random}};
    uw_array = {1{$random}};
    sw_array = {1{$random}};
    ur_array = {1{$random}};
    sr_array = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
`endif

  assign T32 = T2 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T155 : T33;
  assign T33 = T34[1'h1:1'h0];
  assign T34 = {T57, T35};
  assign T35 = T40 & T36;
  assign T36 = T37 - 1'h1;
  assign T37 = 1'h1 << T38;
  assign T38 = T39 + 2'h1;
  assign T39 = T57 - T57;
  assign T40 = R41 >> T57;
  assign T42 = T56 ? T43 : R41;
  assign T43 = T51 | T44;
  assign T44 = T50 ? 4'h0 : T45;
  assign T45 = T46[2'h3:1'h0];
  assign T46 = 4'h1 << T47;
  assign T47 = {1'h1, T48};
  assign T48 = T149[1'h1:1'h1];
  assign T149 = {T154, T150};
  assign T150 = T151[1'h1:1'h1];
  assign T151 = T153 | T152;
  assign T152 = tag_cam_io_hits[1'h1:1'h0];
  assign T153 = tag_cam_io_hits[2'h3:2'h2];
  assign T154 = T153 != 2'h0;
  assign T50 = T149[1'h0:1'h0];
  assign T51 = T53 & T52;
  assign T52 = ~ T45;
  assign T53 = T55 | T54;
  assign T54 = T48 ? 4'h0 : 4'h2;
  assign T55 = R41 & 4'hd;
  assign T56 = io_req_valid & tlb_hit;
  assign tlb_hit = io_ptw_status_vm & tag_cam_io_hit;
  assign T57 = {1'h1, T58};
  assign T58 = R41[1'h1:1'h1];
  assign T155 = T160 ? 1'h0 : T156;
  assign T156 = T159 ? 1'h1 : T157;
  assign T157 = T158 ? 2'h2 : 2'h3;
  assign T158 = T59[2'h2:2'h2];
  assign T59 = ~ tag_cam_io_valid_bits;
  assign T159 = T59[1'h1:1'h1];
  assign T160 = T59[1'h0:1'h0];
  assign has_invalid_entry = T60 ^ 1'h1;
  assign T60 = tag_cam_io_valid_bits == 4'hf;
  assign T2 = T8 & tlb_miss;
  assign tlb_miss = T6 & T3;
  assign T3 = bad_va ^ 1'h1;
  assign bad_va = T5 != T4;
  assign T4 = io_req_bits_vpn[5'h1d:5'h1d];
  assign T5 = io_req_bits_vpn[5'h1e:5'h1e];
  assign T6 = io_ptw_status_vm & T7;
  assign T7 = tag_cam_io_hit ^ 1'h1;
  assign T8 = io_req_ready & io_req_valid;
  assign T168 = r_refill_tag[6'h24:1'h0];
  assign T0 = T2 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T1;
  assign T1 = {io_req_bits_asid, io_req_bits_vpn};
  assign T169 = T170 & io_ptw_resp_valid;
  assign T170 = state == 2'h2;
  assign T148 = reset ? 2'h0 : T10;
  assign T10 = io_ptw_resp_valid ? 2'h0 : T11;
  assign T11 = T20 ? 2'h3 : T12;
  assign T12 = T19 ? 2'h3 : T13;
  assign T13 = T18 ? 2'h2 : T14;
  assign T14 = T16 ? 2'h0 : T15;
  assign T15 = T2 ? 2'h1 : state;
  assign T16 = T17 & io_ptw_invalidate;
  assign T17 = state == 2'h1;
  assign T18 = T17 & io_ptw_req_ready;
  assign T19 = T18 & io_ptw_invalidate;
  assign T20 = T21 & io_ptw_invalidate;
  assign T21 = state == 2'h2;
  assign T171 = lookup_tag[6'h24:1'h0];
  assign T172 = T175 & T173;
  assign T173 = io_req_bits_instruction ? io_resp_xcpt_if : T174;
  assign T174 = io_resp_xcpt_ld & io_resp_xcpt_st;
  assign T175 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits = T147;
  assign T147 = r_refill_tag[5'h1d:1'h0];
  assign io_ptw_req_valid = T9;
  assign T9 = state == 2'h1;
  assign io_resp_xcpt_if = T22;
  assign T22 = bad_va | T23;
  assign T23 = tlb_hit & T24;
  assign T24 = T25 ^ 1'h1;
  assign T25 = io_ptw_status_s ? T68 : T26;
  assign T26 = T27 != 4'h0;
  assign T27 = ux_array & tag_cam_io_hits;
  assign T28 = io_ptw_resp_valid ? T29 : ux_array;
  assign T29 = T66 | T30;
  assign T30 = T161 & T31;
  assign T31 = 1'h1 << r_refill_waddr;
  assign T161 = T61 ? 4'hf : 4'h0;
  assign T61 = T62;
  assign T62 = T63[2'h2:2'h2];
  assign T63 = T162 & io_ptw_resp_bits_perm;
  assign T162 = T64 ? 6'h3f : 6'h0;
  assign T64 = T65;
  assign T65 = io_ptw_resp_bits_error ^ 1'h1;
  assign T66 = ux_array & T67;
  assign T67 = ~ T31;
  assign T68 = T69 != 4'h0;
  assign T69 = sx_array & tag_cam_io_hits;
  assign T70 = io_ptw_resp_valid ? T71 : sx_array;
  assign T71 = T76 | T72;
  assign T72 = T163 & T73;
  assign T73 = 1'h1 << r_refill_waddr;
  assign T163 = T74 ? 4'hf : 4'h0;
  assign T74 = T75;
  assign T75 = T63[3'h5:3'h5];
  assign T76 = sx_array & T77;
  assign T77 = ~ T73;
  assign io_resp_xcpt_st = T78;
  assign T78 = bad_va | T79;
  assign T79 = tlb_hit & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = io_ptw_status_s ? T92 : T82;
  assign T82 = T83 != 4'h0;
  assign T83 = uw_array & tag_cam_io_hits;
  assign T84 = io_ptw_resp_valid ? T85 : uw_array;
  assign T85 = T90 | T86;
  assign T86 = T164 & T87;
  assign T87 = 1'h1 << r_refill_waddr;
  assign T164 = T88 ? 4'hf : 4'h0;
  assign T88 = T89;
  assign T89 = T63[1'h1:1'h1];
  assign T90 = uw_array & T91;
  assign T91 = ~ T87;
  assign T92 = T93 != 4'h0;
  assign T93 = sw_array & tag_cam_io_hits;
  assign T94 = io_ptw_resp_valid ? T95 : sw_array;
  assign T95 = T100 | T96;
  assign T96 = T165 & T97;
  assign T97 = 1'h1 << r_refill_waddr;
  assign T165 = T98 ? 4'hf : 4'h0;
  assign T98 = T99;
  assign T99 = T63[3'h4:3'h4];
  assign T100 = sw_array & T101;
  assign T101 = ~ T97;
  assign io_resp_xcpt_ld = T102;
  assign T102 = bad_va | T103;
  assign T103 = tlb_hit & T104;
  assign T104 = T105 ^ 1'h1;
  assign T105 = io_ptw_status_s ? T116 : T106;
  assign T106 = T107 != 4'h0;
  assign T107 = ur_array & tag_cam_io_hits;
  assign T108 = io_ptw_resp_valid ? T109 : ur_array;
  assign T109 = T114 | T110;
  assign T110 = T166 & T111;
  assign T111 = 1'h1 << r_refill_waddr;
  assign T166 = T112 ? 4'hf : 4'h0;
  assign T112 = T113;
  assign T113 = T63[1'h0:1'h0];
  assign T114 = ur_array & T115;
  assign T115 = ~ T111;
  assign T116 = T117 != 4'h0;
  assign T117 = sr_array & tag_cam_io_hits;
  assign T118 = io_ptw_resp_valid ? T119 : sr_array;
  assign T119 = T124 | T120;
  assign T120 = T167 & T121;
  assign T121 = 1'h1 << r_refill_waddr;
  assign T167 = T122 ? 4'hf : 4'h0;
  assign T122 = T123;
  assign T123 = T63[2'h3:2'h3];
  assign T124 = sr_array & T125;
  assign T125 = ~ T121;
  assign io_resp_ppn = T126;
  assign T126 = T144 ? T128 : T127;
  assign T127 = io_req_bits_vpn[5'h12:1'h0];
  assign T128 = T133 | T129;
  assign T129 = T132 ? T130 : 19'h0;
  assign T130 = tag_ram[2'h3];
  assign T132 = tag_cam_io_hits[2'h3:2'h3];
  assign T133 = T137 | T134;
  assign T134 = T136 ? T135 : 19'h0;
  assign T135 = tag_ram[2'h2];
  assign T136 = tag_cam_io_hits[2'h2:2'h2];
  assign T137 = T141 | T138;
  assign T138 = T140 ? T139 : 19'h0;
  assign T139 = tag_ram[2'h1];
  assign T140 = tag_cam_io_hits[1'h1:1'h1];
  assign T141 = T143 ? T142 : 19'h0;
  assign T142 = tag_ram[2'h0];
  assign T143 = tag_cam_io_hits[1'h0:1'h0];
  assign T144 = io_ptw_status_vm & T145;
  assign T145 = io_req_bits_passthrough ^ 1'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T146;
  assign T146 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( io_ptw_invalidate ),
       .io_clear_hit( T172 ),
       .io_tag( T171 ),
       .io_hit( tag_cam_io_hit ),
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T169 ),
       .io_write_tag( T168 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T2) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T56) begin
      R41 <= T43;
    end
    if(T2) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T20) begin
      state <= 2'h3;
    end else if(T19) begin
      state <= 2'h3;
    end else if(T18) begin
      state <= 2'h2;
    end else if(T16) begin
      state <= 2'h0;
    end else if(T2) begin
      state <= 2'h1;
    end
    if(io_ptw_resp_valid) begin
      ux_array <= T29;
    end
    if(io_ptw_resp_valid) begin
      sx_array <= T71;
    end
    if(io_ptw_resp_valid) begin
      uw_array <= T85;
    end
    if(io_ptw_resp_valid) begin
      sw_array <= T95;
    end
    if(io_ptw_resp_valid) begin
      ur_array <= T109;
    end
    if(io_ptw_resp_valid) begin
      sr_array <= T119;
    end
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_ppn;
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [43:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[43:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_xcpt_ma,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output[42:0] io_cpu_btb_resp_bits_target,
    output[2:0] io_cpu_btb_resp_bits_entry,
    output[3:0] io_cpu_btb_resp_bits_bht_index,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input [42:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [2:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [3:0] io_cpu_btb_update_bits_prediction_bits_bht_index,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [42:0] io_cpu_btb_update_bits_pc,
    input [42:0] io_cpu_btb_update_bits_target,
    input [42:0] io_cpu_btb_update_bits_returnAddr,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isCall,
    input  io_cpu_btb_update_bits_isReturn,
    input  io_cpu_btb_update_bits_incorrectTarget,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    input  io_cpu_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id
);

  wire[30:0] T38;
  wire[43:0] s1_pc;
  reg [43:0] s1_pc_;
  wire[43:0] T19;
  wire[43:0] T20;
  wire[43:0] npc;
  wire[43:0] T21;
  wire[43:0] predicted_npc;
  wire[43:0] pcp4;
  wire[42:0] T22;
  wire[43:0] pcp4_0;
  wire T23;
  wire T24;
  wire T25;
  wire[43:0] btbTarget;
  wire T26;
  reg [43:0] s2_pc;
  wire[43:0] T36;
  wire[43:0] T18;
  wire T2;
  wire T3;
  wire icmiss;
  wire T4;
  reg  s2_valid;
  wire T33;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire stall;
  wire T9;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  reg  s1_same_block;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire s0_same_block;
  wire T48;
  wire[43:0] T49;
  wire[43:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[12:0] T59;
  wire[43:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire[42:0] T65;
  wire[43:0] T66;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T0;
  wire T1;
  reg [3:0] s2_btb_resp_bits_bht_index;
  wire[3:0] T10;
  reg [2:0] s2_btb_resp_bits_entry;
  wire[2:0] T11;
  reg [42:0] s2_btb_resp_bits_target;
  wire[42:0] T12;
  reg  s2_btb_resp_bits_taken;
  wire T13;
  reg  s2_btb_resp_valid;
  wire T34;
  wire T14;
  reg  s2_xcpt_if;
  wire T35;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire[31:0] T37;
  wire[127:0] T27;
  wire[6:0] T28;
  wire[1:0] T29;
  wire[43:0] T30;
  wire T31;
  wire T32;
  wire btb_io_resp_valid;
  wire btb_io_resp_bits_taken;
  wire[42:0] btb_io_resp_bits_target;
  wire[2:0] btb_io_resp_bits_entry;
  wire[3:0] btb_io_resp_bits_bht_index;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire icache_io_resp_valid;
  wire[127:0] icache_io_resp_bits_datablock;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire[1:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire[2:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[5:0] icache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] icache_io_mem_acquire_bits_payload_subword_addr;
  wire[3:0] icache_io_mem_acquire_bits_payload_atomic_opcode;
  wire icache_io_mem_grant_ready;
  wire icache_io_mem_finish_valid;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[2:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire tlb_io_resp_miss;
  wire[18:0] tlb_io_resp_ppn;
  wire tlb_io_resp_xcpt_if;
  wire tlb_io_ptw_req_valid;
  wire[29:0] tlb_io_ptw_req_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s1_same_block = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_index = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
`endif

  assign T38 = s1_pc >> 4'hd;
  assign s1_pc = s1_pc_ & 44'hffffffffffe;
  assign T19 = io_cpu_req_valid ? io_cpu_req_bits_pc : T20;
  assign T20 = T8 ? npc : s1_pc_;
  assign npc = T21;
  assign T21 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : pcp4;
  assign pcp4 = {T23, T22};
  assign T22 = pcp4_0[6'h2a:1'h0];
  assign pcp4_0 = s1_pc + 44'h4;
  assign T23 = T25 & T24;
  assign T24 = pcp4_0[6'h2a:6'h2a];
  assign T25 = s1_pc[6'h2a:6'h2a];
  assign btbTarget = {T26, btb_io_resp_bits_target};
  assign T26 = btb_io_resp_bits_target[6'h2a:6'h2a];
  assign T36 = reset ? 44'h2000 : T18;
  assign T18 = T2 ? s1_pc : s2_pc;
  assign T2 = T8 & T3;
  assign T3 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T4;
  assign T4 = icache_io_resp_valid ^ 1'h1;
  assign T33 = reset ? 1'h1 : T5;
  assign T5 = io_cpu_req_valid ? 1'h0 : T6;
  assign T6 = T8 ? T7 : s2_valid;
  assign T7 = icmiss ^ 1'h1;
  assign T8 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T9;
  assign T9 = io_cpu_resp_ready ^ 1'h1;
  assign T39 = T41 & T40;
  assign T40 = icmiss ^ 1'h1;
  assign T41 = stall ^ 1'h1;
  assign T42 = T56 & T43;
  assign T43 = s1_same_block ^ 1'h1;
  assign T44 = io_cpu_req_valid ? 1'h0 : T45;
  assign T45 = T8 ? T46 : s1_same_block;
  assign T46 = s0_same_block & T47;
  assign T47 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T51 & T48;
  assign T48 = T50 == T49;
  assign T49 = s1_pc & 44'h10;
  assign T50 = pcp4 & 44'h10;
  assign T51 = T53 & T52;
  assign T52 = btb_io_resp_bits_taken ^ 1'h1;
  assign T53 = T55 & T54;
  assign T54 = io_cpu_req_valid ^ 1'h1;
  assign T55 = icmiss ^ 1'h1;
  assign T56 = stall ^ 1'h1;
  assign T57 = T58 | icmiss;
  assign T58 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T59 = T60[4'hc:1'h0];
  assign T60 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign T61 = T63 & T62;
  assign T62 = s0_same_block ^ 1'h1;
  assign T63 = stall ^ 1'h1;
  assign T64 = io_cpu_invalidate | io_cpu_ptw_invalidate;
  assign T65 = T66[6'h2a:1'h0];
  assign T66 = s1_pc & 44'hffffffffffc;
  assign io_mem_finish_bits_payload_master_xact_id = icache_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = icache_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = icache_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = icache_io_mem_finish_valid;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = icache_io_mem_acquire_bits_payload_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = icache_io_mem_acquire_bits_payload_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = icache_io_mem_acquire_bits_payload_write_mask;
  assign io_mem_acquire_bits_payload_a_type = icache_io_mem_acquire_bits_payload_a_type;
  assign io_mem_acquire_bits_payload_data = icache_io_mem_acquire_bits_payload_data;
  assign io_mem_acquire_bits_payload_client_xact_id = icache_io_mem_acquire_bits_payload_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = icache_io_mem_acquire_bits_payload_addr;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_cpu_ptw_req_bits = tlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T0 = T1 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T1 = T2 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_index = s2_btb_resp_bits_bht_index;
  assign T10 = T1 ? btb_io_resp_bits_bht_index : s2_btb_resp_bits_bht_index;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T11 = T1 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T12 = T1 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T13 = T1 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T34 = reset ? 1'h0 : T14;
  assign T14 = T2 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T35 = reset ? 1'h0 : T15;
  assign T15 = T2 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_xcpt_ma = T16;
  assign T16 = T17 != 2'h0;
  assign T17 = s2_pc[1'h1:1'h0];
  assign io_cpu_resp_bits_data = T37;
  assign T37 = T27[5'h1f:1'h0];
  assign T27 = icache_io_resp_bits_datablock >> T28;
  assign T28 = T29 << 3'h5;
  assign T29 = s2_pc[2'h3:2'h2];
  assign io_cpu_resp_bits_pc = T30;
  assign T30 = s2_pc & 44'hffffffffffc;
  assign io_cpu_resp_valid = T31;
  assign T31 = s2_valid & T32;
  assign T32 = s2_xcpt_if | icache_io_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req( T65 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_index( btb_io_resp_bits_bht_index ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_update_valid( io_cpu_btb_update_valid ),
       .io_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_update_bits_prediction_bits_bht_index( io_cpu_btb_update_bits_prediction_bits_bht_index ),
       .io_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_update_bits_returnAddr( io_cpu_btb_update_bits_returnAddr ),
       .io_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_update_bits_isCall( io_cpu_btb_update_bits_isCall ),
       .io_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_update_bits_incorrectTarget( io_cpu_btb_update_bits_incorrectTarget ),
       .io_invalidate( T64 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T61 ),
       .io_req_bits_idx( T59 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T57 ),
       .io_resp_ready( T42 ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T39 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T38 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_resp_miss( tlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits( tlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T8) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 44'h2000;
    end else if(T2) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T8) begin
      s2_valid <= T7;
    end
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T8) begin
      s1_same_block <= T46;
    end
    if(T1) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T1) begin
      s2_btb_resp_bits_bht_index <= btb_io_resp_bits_bht_index;
    end
    if(T1) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T1) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T1) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T2) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T2) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [19:0] io_req_bits_tag,
    input [5:0] io_req_bits_idx,
    input  io_req_bits_way_en,
    input [1:0] io_req_bits_client_xact_id,
    input [2:0] io_req_bits_master_xact_id,
    input [2:0] io_req_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output io_data_req_bits_way_en,
    output[11:0] io_data_req_bits_addr,
    input [127:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[25:0] io_release_bits_addr,
    output[1:0] io_release_bits_client_xact_id,
    output[2:0] io_release_bits_master_xact_id,
    output[511:0] io_release_bits_data,
    output[2:0] io_release_bits_r_type
);

  reg [2:0] req_r_type;
  wire[2:0] T0;
  wire T1;
  reg [511:0] R2;
  wire[511:0] T3;
  wire[511:0] T4;
  wire[383:0] T5;
  wire T6;
  reg  r2_data_req_fired;
  wire T38;
  wire T7;
  reg  r1_data_req_fired;
  wire T39;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  reg  active;
  wire T40;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [2:0] cnt;
  wire[2:0] T41;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  reg [2:0] req_master_xact_id;
  wire[2:0] T26;
  reg [1:0] req_client_xact_id;
  wire[1:0] T27;
  wire[25:0] T28;
  wire[25:0] T29;
  reg [5:0] req_idx;
  wire[5:0] T30;
  reg [19:0] req_tag;
  wire[19:0] T31;
  wire[11:0] T32;
  wire[7:0] T33;
  wire[1:0] T34;
  reg  req_way_en;
  wire T35;
  wire fire;
  wire T36;
  wire T37;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_r_type = {1{$random}};
    R2 = {16{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    cnt = {1{$random}};
    req_master_xact_id = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_idx = {1{$random}};
    req_tag = {1{$random}};
    req_way_en = {1{$random}};
  end
`endif

  assign io_release_bits_r_type = req_r_type;
  assign T0 = T1 ? io_req_bits_r_type : req_r_type;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_data = R2;
  assign T3 = T6 ? T4 : R2;
  assign T4 = {io_data_resp, T5};
  assign T5 = R2[9'h1ff:8'h80];
  assign T6 = active & r2_data_req_fired;
  assign T38 = reset ? 1'h0 : T7;
  assign T7 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T39 = reset ? 1'h0 : T8;
  assign T8 = T10 ? 1'h1 : T9;
  assign T9 = active ? 1'h0 : r1_data_req_fired;
  assign T10 = active & T11;
  assign T11 = T13 & T12;
  assign T12 = io_meta_read_ready & io_meta_read_valid;
  assign T13 = io_data_req_ready & io_data_req_valid;
  assign T40 = reset ? 1'h0 : T14;
  assign T14 = T1 ? 1'h1 : T15;
  assign T15 = T17 ? T16 : active;
  assign T16 = io_release_ready ^ 1'h1;
  assign T17 = active & T18;
  assign T18 = T23 & T19;
  assign T19 = cnt == 3'h4;
  assign T41 = reset ? 3'h0 : T20;
  assign T20 = T1 ? 3'h0 : T21;
  assign T21 = T10 ? T22 : cnt;
  assign T22 = cnt + 3'h1;
  assign T23 = T25 & T24;
  assign T24 = r2_data_req_fired ^ 1'h1;
  assign T25 = r1_data_req_fired ^ 1'h1;
  assign io_release_bits_master_xact_id = req_master_xact_id;
  assign T26 = T1 ? io_req_bits_master_xact_id : req_master_xact_id;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T27 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr = T28;
  assign T28 = T29;
  assign T29 = {req_tag, req_idx};
  assign T30 = T1 ? io_req_bits_idx : req_idx;
  assign T31 = T1 ? io_req_bits_tag : req_tag;
  assign io_release_valid = T17;
  assign io_data_req_bits_addr = T32;
  assign T32 = T33 << 3'h4;
  assign T33 = {req_idx, T34};
  assign T34 = cnt[1'h1:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T35 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T36;
  assign T36 = cnt < 3'h4;
  assign io_meta_read_bits_tag = req_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T37;
  assign T37 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(T6) begin
      R2 <= T4;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T10) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T17) begin
      active <= T16;
    end
    if(reset) begin
      cnt <= 3'h0;
    end else if(T1) begin
      cnt <= 3'h0;
    end else if(T10) begin
      cnt <= T22;
    end
    if(T1) begin
      req_master_xact_id <= io_req_bits_master_xact_id;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_idx <= io_req_bits_idx;
    end
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr,
    input [2:0] io_req_bits_master_xact_id,
    input [1:0] io_req_bits_p_type,
    input [1:0] io_req_bits_client_xact_id,
    input  io_rep_ready,
    output io_rep_valid,
    output[25:0] io_rep_bits_addr,
    output[1:0] io_rep_bits_client_xact_id,
    output[2:0] io_rep_bits_master_xact_id,
    output[511:0] io_rep_bits_data,
    output[2:0] io_rep_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    input  io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_line_state_state
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  reg [1:0] req_p_type;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg [3:0] state;
  wire[3:0] T93;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] T27;
  wire T28;
  reg [1:0] line_state_state;
  wire[1:0] T29;
  wire T30;
  wire hit;
  reg  way_en;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire[2:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  wire[1:0] T49;
  reg [2:0] req_master_xact_id;
  wire[2:0] T50;
  reg [1:0] req_client_xact_id;
  wire[1:0] T51;
  wire[5:0] T94;
  reg [25:0] req_addr;
  wire[25:0] T52;
  wire[19:0] T53;
  wire T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[19:0] T62;
  wire[5:0] T95;
  wire T63;
  wire[19:0] T64;
  wire[5:0] T96;
  wire T65;
  wire[2:0] T66;
  wire[2:0] T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire[2:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire[2:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire[511:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[25:0] T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_p_type = {1{$random}};
    state = {1{$random}};
    line_state_state = {1{$random}};
    way_en = {1{$random}};
    req_master_xact_id = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr = {1{$random}};
  end
`endif

  assign io_wb_req_bits_r_type = T0;
  assign T0 = T47 ? T41 : T1;
  assign T1 = T40 ? 3'h4 : T2;
  assign T2 = T39 ? 3'h5 : T3;
  assign T3 = T4 ? 3'h6 : 3'h4;
  assign T4 = req_p_type == 2'h2;
  assign T5 = T6 ? io_req_bits_p_type : req_p_type;
  assign T6 = T7 & io_req_valid;
  assign T7 = state == 4'h1;
  assign T93 = reset ? 4'h1 : T8;
  assign T8 = T38 ? 4'h1 : T9;
  assign T9 = T6 ? 4'h2 : T10;
  assign T10 = T36 ? 4'h3 : T11;
  assign T11 = T35 ? 4'h4 : T12;
  assign T12 = T33 ? 4'h2 : T13;
  assign T13 = T32 ? 4'h5 : T14;
  assign T14 = T30 ? T27 : T15;
  assign T15 = T25 ? 4'h1 : T16;
  assign T16 = T23 ? 4'h7 : T17;
  assign T17 = T21 ? 4'h8 : T18;
  assign T18 = T19 ? 4'h1 : state;
  assign T19 = T20 & io_meta_write_ready;
  assign T20 = state == 4'h8;
  assign T21 = T22 & io_wb_req_ready;
  assign T22 = state == 4'h7;
  assign T23 = T24 & io_wb_req_ready;
  assign T24 = state == 4'h6;
  assign T25 = T26 & io_rep_ready;
  assign T26 = state == 4'h5;
  assign T27 = T28 ? 4'h6 : 4'h8;
  assign T28 = line_state_state == 2'h3;
  assign T29 = T32 ? io_line_state_state : line_state_state;
  assign T30 = T25 & hit;
  assign hit = way_en != 1'h0;
  assign T31 = T32 ? io_way_en : way_en;
  assign T32 = state == 4'h4;
  assign T33 = T32 & T34;
  assign T34 = io_mshr_rdy ^ 1'h1;
  assign T35 = state == 4'h3;
  assign T36 = T37 & io_meta_read_ready;
  assign T37 = state == 4'h2;
  assign T38 = state == 4'h0;
  assign T39 = req_p_type == 2'h1;
  assign T40 = req_p_type == 2'h0;
  assign T41 = T46 ? 3'h1 : T42;
  assign T42 = T45 ? 3'h2 : T43;
  assign T43 = T44 ? 3'h3 : 3'h1;
  assign T44 = req_p_type == 2'h2;
  assign T45 = req_p_type == 2'h1;
  assign T46 = req_p_type == 2'h0;
  assign T47 = T48 == 2'h3;
  assign T48 = hit ? line_state_state : T49;
  assign T49 = 2'h0;
  assign io_wb_req_bits_master_xact_id = req_master_xact_id;
  assign T50 = T6 ? io_req_bits_master_xact_id : req_master_xact_id;
  assign io_wb_req_bits_client_xact_id = req_client_xact_id;
  assign T51 = T6 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_wb_req_bits_way_en = way_en;
  assign io_wb_req_bits_idx = T94;
  assign T94 = req_addr[3'h5:1'h0];
  assign T52 = T6 ? io_req_bits_addr : req_addr;
  assign io_wb_req_bits_tag = T53;
  assign T53 = req_addr >> 3'h6;
  assign io_wb_req_valid = T54;
  assign T54 = state == 4'h6;
  assign io_meta_write_bits_data_coh_state = T55;
  assign T55 = T56;
  assign T56 = T61 ? 2'h0 : T57;
  assign T57 = T60 ? 2'h1 : T58;
  assign T58 = T59 ? line_state_state : line_state_state;
  assign T59 = req_p_type == 2'h2;
  assign T60 = req_p_type == 2'h1;
  assign T61 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T62;
  assign T62 = req_addr >> 3'h6;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T95;
  assign T95 = req_addr[3'h5:1'h0];
  assign io_meta_write_valid = T63;
  assign T63 = state == 4'h8;
  assign io_meta_read_bits_tag = T64;
  assign T64 = req_addr >> 3'h6;
  assign io_meta_read_bits_idx = T96;
  assign T96 = req_addr[3'h5:1'h0];
  assign io_meta_read_valid = T65;
  assign T65 = state == 4'h2;
  assign io_rep_bits_r_type = T66;
  assign T66 = T67;
  assign T67 = T80 ? T74 : T68;
  assign T68 = T73 ? 3'h4 : T69;
  assign T69 = T72 ? 3'h5 : T70;
  assign T70 = T71 ? 3'h6 : 3'h4;
  assign T71 = req_p_type == 2'h2;
  assign T72 = req_p_type == 2'h1;
  assign T73 = req_p_type == 2'h0;
  assign T74 = T79 ? 3'h1 : T75;
  assign T75 = T78 ? 3'h2 : T76;
  assign T76 = T77 ? 3'h3 : 3'h1;
  assign T77 = req_p_type == 2'h2;
  assign T78 = req_p_type == 2'h1;
  assign T79 = req_p_type == 2'h0;
  assign T80 = T81 == 2'h3;
  assign T81 = hit ? line_state_state : T82;
  assign T82 = 2'h0;
  assign io_rep_bits_data = T83;
  assign T83 = 512'h0;
  assign io_rep_bits_master_xact_id = T84;
  assign T84 = req_master_xact_id;
  assign io_rep_bits_client_xact_id = T85;
  assign T85 = req_client_xact_id;
  assign io_rep_bits_addr = T86;
  assign T86 = req_addr;
  assign io_rep_valid = T87;
  assign T87 = T91 & T88;
  assign T88 = T89 ^ 1'h1;
  assign T89 = hit & T90;
  assign T90 = line_state_state == 2'h3;
  assign T91 = state == 4'h5;
  assign io_req_ready = T92;
  assign T92 = state == 4'h1;

  always @(posedge clk) begin
    if(T6) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(reset) begin
      state <= 4'h1;
    end else if(T38) begin
      state <= 4'h1;
    end else if(T6) begin
      state <= 4'h2;
    end else if(T36) begin
      state <= 4'h3;
    end else if(T35) begin
      state <= 4'h4;
    end else if(T33) begin
      state <= 4'h2;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T30) begin
      state <= T27;
    end else if(T25) begin
      state <= 4'h1;
    end else if(T23) begin
      state <= 4'h7;
    end else if(T21) begin
      state <= 4'h8;
    end else if(T19) begin
      state <= 4'h1;
    end
    if(T32) begin
      line_state_state <= io_line_state_state;
    end
    if(T32) begin
      way_en <= io_way_en;
    end
    if(T6) begin
      req_master_xact_id <= io_req_bits_master_xact_id;
    end
    if(T6) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T6) begin
      req_addr <= io_req_bits_addr;
    end
  end
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [19:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [19:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[19:0] io_out_bits_tag,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[19:0] T2;
  wire T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T2;
  assign T2 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T3 = T0;
  assign io_out_bits_idx = T4;
  assign T4 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input  io_in_1_bits_way_en,
    input [19:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_in_0_bits_way_en,
    input [19:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output io_out_bits_way_en,
    output[19:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[1:0] T2;
  wire T3;
  wire[19:0] T4;
  wire T5;
  wire[5:0] T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T2;
  assign T2 = T3 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T3 = T0;
  assign io_out_bits_data_tag = T4;
  assign T4 = T3 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T5;
  assign T5 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T6;
  assign T6 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_7(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_client_xact_id,
    input [511:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_a_type,
    input [5:0] io_in_1_bits_write_mask,
    input [2:0] io_in_1_bits_subword_addr,
    input [3:0] io_in_1_bits_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_client_xact_id,
    input [511:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_a_type,
    input [5:0] io_in_0_bits_write_mask,
    input [2:0] io_in_0_bits_subword_addr,
    input [3:0] io_in_0_bits_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[1:0] io_out_bits_client_xact_id,
    output[511:0] io_out_bits_data,
    output[2:0] io_out_bits_a_type,
    output[5:0] io_out_bits_write_mask,
    output[2:0] io_out_bits_subword_addr,
    output[3:0] io_out_bits_atomic_opcode,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[3:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[5:0] T5;
  wire[2:0] T6;
  wire[511:0] T7;
  wire[1:0] T8;
  wire[25:0] T9;
  wire T10;
  wire T11;
  wire T12;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_atomic_opcode = T2;
  assign T2 = T3 ? io_in_1_bits_atomic_opcode : io_in_0_bits_atomic_opcode;
  assign T3 = T0;
  assign io_out_bits_subword_addr = T4;
  assign T4 = T3 ? io_in_1_bits_subword_addr : io_in_0_bits_subword_addr;
  assign io_out_bits_write_mask = T5;
  assign T5 = T3 ? io_in_1_bits_write_mask : io_in_0_bits_write_mask;
  assign io_out_bits_a_type = T6;
  assign T6 = T3 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_data = T7;
  assign T7 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_client_xact_id = T8;
  assign T8 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T9;
  assign T9 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T10;
  assign T10 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_8(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_payload_master_xact_id = T2;
  assign T2 = T3 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T3 = T0;
  assign io_out_bits_header_dst = T4;
  assign T4 = T3 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T5;
  assign T5 = T3 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T6;
  assign T6 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T7;
  assign T7 = T8 & io_out_ready;
  assign T8 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [19:0] io_in_1_bits_tag,
    input [5:0] io_in_1_bits_idx,
    input  io_in_1_bits_way_en,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_master_xact_id,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [19:0] io_in_0_bits_tag,
    input [5:0] io_in_0_bits_idx,
    input  io_in_0_bits_way_en,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_master_xact_id,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[19:0] io_out_bits_tag,
    output[5:0] io_out_bits_idx,
    output io_out_bits_way_en,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_master_xact_id,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[1:0] T5;
  wire T6;
  wire[5:0] T7;
  wire[19:0] T8;
  wire T9;
  wire T10;
  wire T11;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_master_xact_id = T4;
  assign T4 = T3 ? io_in_1_bits_master_xact_id : io_in_0_bits_master_xact_id;
  assign io_out_bits_client_xact_id = T5;
  assign T5 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_way_en = T6;
  assign T6 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T7;
  assign T7 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_bits_tag = T8;
  assign T8 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_valid = T9;
  assign T9 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_9(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_kill,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_phys,
    input [43:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    input [7:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_kill,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_phys,
    input [43:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input [7:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_kill,
    output[2:0] io_out_bits_typ,
    output io_out_bits_phys,
    output[43:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output[7:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[4:0] T2;
  wire T3;
  wire[4:0] T4;
  wire[7:0] T5;
  wire[63:0] T6;
  wire[43:0] T7;
  wire T8;
  wire[2:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T2;
  assign T2 = T3 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T3 = T0;
  assign io_out_bits_cmd = T4;
  assign T4 = T3 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T5;
  assign T5 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_data = T6;
  assign T6 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_addr = T7;
  assign T7 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_phys = T8;
  assign T8 = T3 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_typ = T9;
  assign T9 = T3 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_kill = T10;
  assign T10 = T3 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_valid = T11;
  assign T11 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T12;
  assign T12 = T13 & io_out_ready;
  assign T13 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_10(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits = T2;
  assign T2 = T3 ? io_in_1_bits : io_in_0_bits;
  assign T3 = T0;
  assign io_out_valid = T4;
  assign T4 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T5;
  assign T5 = T6 & io_out_ready;
  assign T6 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_14(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_kill,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_phys,
    input [43:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input [7:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_kill,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_phys,
    output[43:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data,
    output[7:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T31;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  reg [3:0] R4;
  wire[3:0] T32;
  wire[3:0] T5;
  wire[3:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[4:0] T10;
  wire[130:0] T11;
  reg [130:0] ram [15:0];
  wire[130:0] T12;
  wire[130:0] T13;
  wire[130:0] T14;
  wire[81:0] T15;
  wire[9:0] T16;
  wire[71:0] T17;
  wire[48:0] T18;
  wire[44:0] T19;
  wire[3:0] T20;
  wire[4:0] T21;
  wire[7:0] T22;
  wire[63:0] T23;
  wire[43:0] T24;
  wire T25;
  wire[2:0] T26;
  wire T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 4'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T10;
  assign T10 = T11[3'h4:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_cmd, io_enq_bits_sdq_id};
  assign T17 = {io_enq_bits_data, io_enq_bits_tag};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_phys, io_enq_bits_addr};
  assign T20 = {io_enq_bits_kill, io_enq_bits_typ};
  assign io_deq_bits_cmd = T21;
  assign T21 = T11[4'h9:3'h5];
  assign io_deq_bits_tag = T22;
  assign T22 = T11[5'h11:4'ha];
  assign io_deq_bits_data = T23;
  assign T23 = T11[7'h51:5'h12];
  assign io_deq_bits_addr = T24;
  assign T24 = T11[7'h7d:7'h52];
  assign io_deq_bits_phys = T25;
  assign T25 = T11[7'h7e:7'h7e];
  assign io_deq_bits_typ = T26;
  assign T26 = T11[8'h81:7'h7f];
  assign io_deq_bits_kill = T27;
  assign T27 = T11[8'h82:8'h82];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 4'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    input [4:0] io_req_sdq_id,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    //output[511:0] io_mem_req_bits_data
    output[2:0] io_mem_req_bits_a_type,
    //output[5:0] io_mem_req_bits_write_mask
    //output[2:0] io_mem_req_bits_subword_addr
    //output[3:0] io_mem_req_bits_atomic_opcode
    output io_mem_resp_way_en,
    output[11:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T204;
  wire can_finish;
  wire T81;
  reg [3:0] state;
  wire[3:0] T200;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire refill_done;
  wire T28;
  reg [1:0] refill_count;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire reply;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire T82;
  wire T83;
  wire T84;
  wire T205;
  wire T206;
  wire T207;
  wire wb_done;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T86;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire sec_rdy;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire idx_match;
  wire[5:0] T74;
  wire[5:0] req_idx;
  reg [43:0] req_addr;
  wire[43:0] T75;
  wire T221;
  wire T0;
  wire T1;
  wire T2;
  reg [1:0] meta_hazard;
  wire[1:0] T199;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  reg  req_way_en;
  wire T76;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[4:0] T85;
  wire[43:0] T201;
  wire[31:0] T87;
  wire[31:0] T88;
  wire[11:0] T89;
  wire[5:0] T90;
  wire T91;
  wire T92;
  wire[1:0] T93;
  reg [1:0] line_state_state;
  wire[1:0] T94;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T97;
  wire[1:0] T98;
  wire[1:0] T99;
  wire T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire[1:0] meta_on_flush_state;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire[127:0] T202;
  reg [63:0] req_data;
  wire[63:0] T118;
  wire[11:0] T119;
  wire[7:0] T120;
  reg [2:0] acquire_type;
  wire[2:0] T121;
  wire[2:0] T122;
  wire[2:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[2:0] T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[25:0] T148;
  wire[25:0] T149;
  wire T150;
  wire T151;
  wire[19:0] T203;
  wire[31:0] T152;
  wire T153;
  wire T154;
  wire T155;
  wire T198;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire rpq_io_deq_bits_kill;
  wire[2:0] rpq_io_deq_bits_typ;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[63:0] rpq_io_deq_bits_data;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire ackq_io_enq_ready;
  wire ackq_io_deq_valid;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[2:0] ackq_io_deq_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    req_data = {2{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T204 = io_mem_finish_ready & can_finish;
  assign can_finish = T82 | T81;
  assign T81 = state == 4'h5;
  assign T200 = reset ? 4'h0 : T10;
  assign T10 = T68 ? T66 : T11;
  assign T11 = T64 ? 4'h4 : T12;
  assign T12 = T42 ? 4'h6 : T13;
  assign T13 = T41 ? 4'h2 : T14;
  assign T14 = T39 ? 4'h3 : T15;
  assign T15 = T37 ? 4'h4 : T16;
  assign T16 = T36 ? 4'h5 : T17;
  assign T17 = T27 ? 4'h6 : T18;
  assign T18 = T25 ? 4'h7 : T19;
  assign T19 = T24 ? 4'h8 : T20;
  assign T20 = T21 ? 4'h0 : state;
  assign T21 = T23 & T22;
  assign T22 = rpq_io_deq_valid ^ 1'h1;
  assign T23 = state == 4'h8;
  assign T24 = state == 4'h7;
  assign T25 = T26 & io_meta_write_ready;
  assign T26 = state == 4'h6;
  assign T27 = T35 & refill_done;
  assign refill_done = reply & T28;
  assign T28 = refill_count == 2'h3;
  assign T29 = T33 ? 2'h0 : T30;
  assign T30 = T32 ? T31 : refill_count;
  assign T31 = refill_count + 2'h1;
  assign T32 = T35 & reply;
  assign T33 = io_req_pri_val & io_req_pri_rdy;
  assign reply = io_mem_grant_valid & T34;
  assign T34 = io_mem_grant_bits_payload_client_xact_id == 2'h0;
  assign T35 = state == 4'h5;
  assign T36 = io_mem_req_ready & io_mem_req_valid;
  assign T37 = T38 & io_meta_write_ready;
  assign T38 = state == 4'h3;
  assign T39 = T40 & reply;
  assign T40 = state == 4'h2;
  assign T41 = io_wb_req_ready & io_wb_req_valid;
  assign T42 = T63 & T43;
  assign T43 = T52 ? T49 : T44;
  assign T44 = T46 | T45;
  assign T45 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T46 = T48 | T47;
  assign T47 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T48 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T49 = T51 | T50;
  assign T50 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T51 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T52 = T54 | T53;
  assign T53 = io_req_bits_cmd == 5'h6;
  assign T54 = T56 | T55;
  assign T55 = io_req_bits_cmd == 5'h3;
  assign T56 = T60 | T57;
  assign T57 = T59 | T58;
  assign T58 = io_req_bits_cmd == 5'h4;
  assign T59 = io_req_bits_cmd[2'h3:2'h3];
  assign T60 = T62 | T61;
  assign T61 = io_req_bits_cmd == 5'h7;
  assign T62 = io_req_bits_cmd == 5'h1;
  assign T63 = T33 & io_req_bits_tag_match;
  assign T64 = T63 & T65;
  assign T65 = T43 ^ 1'h1;
  assign T66 = T67 ? 4'h1 : 4'h3;
  assign T67 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T68 = T33 & T69;
  assign T69 = io_req_bits_tag_match ^ 1'h1;
  assign T82 = T84 | T83;
  assign T83 = state == 4'h4;
  assign T84 = state == 4'h0;
  assign T205 = T207 & T206;
  assign T206 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T207 = wb_done | refill_done;
  assign wb_done = reply & T208;
  assign T208 = state == 4'h2;
  assign T209 = T86 ? 1'h0 : T210;
  assign T210 = T212 | T211;
  assign T211 = state == 4'h0;
  assign T212 = io_replay_ready & T213;
  assign T213 = state == 4'h8;
  assign T86 = io_meta_read_ready ^ 1'h1;
  assign T214 = T219 & T215;
  assign T215 = T216 ^ 1'h1;
  assign T216 = T218 | T217;
  assign T217 = io_req_bits_cmd == 5'h3;
  assign T218 = io_req_bits_cmd == 5'h2;
  assign T219 = T221 | T220;
  assign T220 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T156;
  assign T156 = T193 | T157;
  assign T157 = T190 & T158;
  assign T158 = T159 ^ 1'h1;
  assign T159 = T173 | T160;
  assign T160 = T162 & T161;
  assign T161 = io_mem_req_bits_a_type != 3'h1;
  assign T162 = T164 | T163;
  assign T163 = io_req_bits_cmd == 5'h6;
  assign T164 = T166 | T165;
  assign T165 = io_req_bits_cmd == 5'h3;
  assign T166 = T170 | T167;
  assign T167 = T169 | T168;
  assign T168 = io_req_bits_cmd == 5'h4;
  assign T169 = io_req_bits_cmd[2'h3:2'h3];
  assign T170 = T172 | T171;
  assign T171 = io_req_bits_cmd == 5'h7;
  assign T172 = io_req_bits_cmd == 5'h1;
  assign T173 = T183 & T174;
  assign T174 = T176 | T175;
  assign T175 = 3'h6 == io_mem_req_bits_a_type;
  assign T176 = T178 | T177;
  assign T177 = 3'h5 == io_mem_req_bits_a_type;
  assign T178 = T180 | T179;
  assign T179 = 3'h4 == io_mem_req_bits_a_type;
  assign T180 = T182 | T181;
  assign T181 = 3'h3 == io_mem_req_bits_a_type;
  assign T182 = 3'h2 == io_mem_req_bits_a_type;
  assign T183 = T187 | T184;
  assign T184 = T186 | T185;
  assign T185 = io_req_bits_cmd == 5'h4;
  assign T186 = io_req_bits_cmd[2'h3:2'h3];
  assign T187 = T189 | T188;
  assign T188 = io_req_bits_cmd == 5'h6;
  assign T189 = io_req_bits_cmd == 5'h0;
  assign T190 = T192 | T191;
  assign T191 = state == 4'h5;
  assign T192 = state == 4'h4;
  assign T193 = T195 | T194;
  assign T194 = state == 4'h3;
  assign T195 = T197 | T196;
  assign T196 = state == 4'h2;
  assign T197 = state == 4'h1;
  assign idx_match = req_idx == T74;
  assign T74 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T75 = T33 ? io_req_bits_addr : req_addr;
  assign T221 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T0;
  assign T0 = T73 | T1;
  assign T1 = T8 & T2;
  assign T2 = meta_hazard == 2'h0;
  assign T199 = reset ? 2'h0 : T3;
  assign T3 = T7 ? 2'h1 : T4;
  assign T4 = T6 ? T5 : meta_hazard;
  assign T5 = meta_hazard + 2'h1;
  assign T6 = meta_hazard != 2'h0;
  assign T7 = io_meta_write_ready & io_meta_write_valid;
  assign T8 = T70 & T9;
  assign T9 = state != 4'h3;
  assign T70 = T72 & T71;
  assign T71 = state != 4'h2;
  assign T72 = state != 4'h1;
  assign T73 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_master_xact_id = 3'h0;
  assign io_wb_req_bits_client_xact_id = 2'h0;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T76 = T33 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = req_idx;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T77 = T33 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T78;
  assign T78 = T79 & ackq_io_enq_ready;
  assign T79 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T80;
  assign T80 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T85;
  assign T85 = T86 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_data = rpq_io_deq_bits_data;
  assign io_replay_bits_addr = T201;
  assign T201 = {12'h0, T87};
  assign T87 = T88;
  assign T88 = {io_tag, T89};
  assign T89 = {req_idx, T90};
  assign T90 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T91;
  assign T91 = T92 & rpq_io_deq_valid;
  assign T92 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T93;
  assign T93 = T113 ? meta_on_flush_state : line_state_state;
  assign T94 = T42 ? meta_on_hit_state : T95;
  assign T95 = T33 ? meta_on_flush_state : T96;
  assign T96 = T32 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T97;
  assign T97 = T104 ? 2'h1 : T98;
  assign T98 = T103 ? T101 : T99;
  assign T99 = T100 ? 2'h3 : 2'h0;
  assign T100 = io_mem_grant_bits_payload_g_type == 4'h5;
  assign T101 = T102 ? 2'h3 : 2'h2;
  assign T102 = io_mem_req_bits_a_type == 3'h1;
  assign T103 = io_mem_grant_bits_payload_g_type == 4'h2;
  assign T104 = io_mem_grant_bits_payload_g_type == 4'h1;
  assign meta_on_hit_state = T105;
  assign T105 = T106 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T106 = T110 | T107;
  assign T107 = T109 | T108;
  assign T108 = io_req_bits_cmd == 5'h4;
  assign T109 = io_req_bits_cmd[2'h3:2'h3];
  assign T110 = T112 | T111;
  assign T111 = io_req_bits_cmd == 5'h7;
  assign T112 = io_req_bits_cmd == 5'h1;
  assign meta_on_flush_state = 2'h0;
  assign T113 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T114;
  assign T114 = T116 | T115;
  assign T115 = state == 4'h3;
  assign T116 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T117;
  assign T117 = state == 4'h8;
  assign io_mem_resp_data = T202;
  assign T202 = {64'h0, req_data};
  assign T118 = T33 ? io_req_bits_data : req_data;
  assign io_mem_resp_addr = T119;
  assign T119 = T120 << 3'h4;
  assign T120 = {req_idx, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_a_type = acquire_type;
  assign T121 = T33 ? T136 : T122;
  assign T122 = T135 ? T123 : acquire_type;
  assign T123 = T124 ? 3'h1 : io_mem_req_bits_a_type;
  assign T124 = T126 | T125;
  assign T125 = io_req_bits_cmd == 5'h6;
  assign T126 = T128 | T127;
  assign T127 = io_req_bits_cmd == 5'h3;
  assign T128 = T132 | T129;
  assign T129 = T131 | T130;
  assign T130 = io_req_bits_cmd == 5'h4;
  assign T131 = io_req_bits_cmd[2'h3:2'h3];
  assign T132 = T134 | T133;
  assign T133 = io_req_bits_cmd == 5'h7;
  assign T134 = io_req_bits_cmd == 5'h1;
  assign T135 = io_req_sec_val & io_req_sec_rdy;
  assign T136 = T137 ? 3'h1 : 3'h0;
  assign T137 = T139 | T138;
  assign T138 = io_req_bits_cmd == 5'h6;
  assign T139 = T141 | T140;
  assign T140 = io_req_bits_cmd == 5'h3;
  assign T141 = T145 | T142;
  assign T142 = T144 | T143;
  assign T143 = io_req_bits_cmd == 5'h4;
  assign T144 = io_req_bits_cmd[2'h3:2'h3];
  assign T145 = T147 | T146;
  assign T146 = io_req_bits_cmd == 5'h7;
  assign T147 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_client_xact_id = 2'h0;
  assign io_mem_req_bits_addr = T148;
  assign T148 = T149;
  assign T149 = {io_tag, req_idx};
  assign io_mem_req_valid = T150;
  assign T150 = T151 & ackq_io_enq_ready;
  assign T151 = state == 4'h4;
  assign io_tag = T203;
  assign T203 = T152[5'h13:1'h0];
  assign T152 = req_addr >> 4'hc;
  assign io_idx_match = T153;
  assign T153 = T154 & idx_match;
  assign T154 = state != 4'h0;
  assign io_req_sec_rdy = T155;
  assign T155 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T198;
  assign T198 = state == 4'h0;
  Queue_14 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T214 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_data( io_req_bits_data ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_sdq_id ),
       .io_deq_ready( T209 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_data( rpq_io_deq_bits_data ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_11 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T205 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T204 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T68) begin
      state <= T66;
    end else if(T64) begin
      state <= 4'h4;
    end else if(T42) begin
      state <= 4'h6;
    end else if(T41) begin
      state <= 4'h2;
    end else if(T39) begin
      state <= 4'h3;
    end else if(T37) begin
      state <= 4'h4;
    end else if(T36) begin
      state <= 4'h5;
    end else if(T27) begin
      state <= 4'h6;
    end else if(T25) begin
      state <= 4'h7;
    end else if(T24) begin
      state <= 4'h8;
    end else if(T21) begin
      state <= 4'h0;
    end
    if(T33) begin
      refill_count <= 2'h0;
    end else if(T32) begin
      refill_count <= T31;
    end
    if(T33) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T7) begin
      meta_hazard <= 2'h1;
    end else if(T6) begin
      meta_hazard <= T5;
    end
    if(T33) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T33) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T42) begin
      line_state_state <= meta_on_hit_state;
    end else if(T33) begin
      line_state_state <= meta_on_flush_state;
    end else if(T32) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T33) begin
      req_data <= io_req_bits_data;
    end
    if(T33) begin
      acquire_type <= T136;
    end else if(T135) begin
      acquire_type <= T123;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    input [4:0] io_req_sdq_id,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    //output[511:0] io_mem_req_bits_data
    output[2:0] io_mem_req_bits_a_type,
    //output[5:0] io_mem_req_bits_write_mask
    //output[2:0] io_mem_req_bits_subword_addr
    //output[3:0] io_mem_req_bits_atomic_opcode
    output io_mem_resp_way_en,
    output[11:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T204;
  wire can_finish;
  wire T81;
  reg [3:0] state;
  wire[3:0] T200;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire refill_done;
  wire T28;
  reg [1:0] refill_count;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire reply;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire T82;
  wire T83;
  wire T84;
  wire T205;
  wire T206;
  wire T207;
  wire wb_done;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T86;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire sec_rdy;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire idx_match;
  wire[5:0] T74;
  wire[5:0] req_idx;
  reg [43:0] req_addr;
  wire[43:0] T75;
  wire T221;
  wire T0;
  wire T1;
  wire T2;
  reg [1:0] meta_hazard;
  wire[1:0] T199;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  reg  req_way_en;
  wire T76;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[4:0] T85;
  wire[43:0] T201;
  wire[31:0] T87;
  wire[31:0] T88;
  wire[11:0] T89;
  wire[5:0] T90;
  wire T91;
  wire T92;
  wire[1:0] T93;
  reg [1:0] line_state_state;
  wire[1:0] T94;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T97;
  wire[1:0] T98;
  wire[1:0] T99;
  wire T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire[1:0] meta_on_flush_state;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire[127:0] T202;
  reg [63:0] req_data;
  wire[63:0] T118;
  wire[11:0] T119;
  wire[7:0] T120;
  reg [2:0] acquire_type;
  wire[2:0] T121;
  wire[2:0] T122;
  wire[2:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[2:0] T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[25:0] T148;
  wire[25:0] T149;
  wire T150;
  wire T151;
  wire[19:0] T203;
  wire[31:0] T152;
  wire T153;
  wire T154;
  wire T155;
  wire T198;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire rpq_io_deq_bits_kill;
  wire[2:0] rpq_io_deq_bits_typ;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[63:0] rpq_io_deq_bits_data;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire ackq_io_enq_ready;
  wire ackq_io_deq_valid;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[2:0] ackq_io_deq_bits_payload_master_xact_id;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    req_data = {2{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T204 = io_mem_finish_ready & can_finish;
  assign can_finish = T82 | T81;
  assign T81 = state == 4'h5;
  assign T200 = reset ? 4'h0 : T10;
  assign T10 = T68 ? T66 : T11;
  assign T11 = T64 ? 4'h4 : T12;
  assign T12 = T42 ? 4'h6 : T13;
  assign T13 = T41 ? 4'h2 : T14;
  assign T14 = T39 ? 4'h3 : T15;
  assign T15 = T37 ? 4'h4 : T16;
  assign T16 = T36 ? 4'h5 : T17;
  assign T17 = T27 ? 4'h6 : T18;
  assign T18 = T25 ? 4'h7 : T19;
  assign T19 = T24 ? 4'h8 : T20;
  assign T20 = T21 ? 4'h0 : state;
  assign T21 = T23 & T22;
  assign T22 = rpq_io_deq_valid ^ 1'h1;
  assign T23 = state == 4'h8;
  assign T24 = state == 4'h7;
  assign T25 = T26 & io_meta_write_ready;
  assign T26 = state == 4'h6;
  assign T27 = T35 & refill_done;
  assign refill_done = reply & T28;
  assign T28 = refill_count == 2'h3;
  assign T29 = T33 ? 2'h0 : T30;
  assign T30 = T32 ? T31 : refill_count;
  assign T31 = refill_count + 2'h1;
  assign T32 = T35 & reply;
  assign T33 = io_req_pri_val & io_req_pri_rdy;
  assign reply = io_mem_grant_valid & T34;
  assign T34 = io_mem_grant_bits_payload_client_xact_id == 2'h1;
  assign T35 = state == 4'h5;
  assign T36 = io_mem_req_ready & io_mem_req_valid;
  assign T37 = T38 & io_meta_write_ready;
  assign T38 = state == 4'h3;
  assign T39 = T40 & reply;
  assign T40 = state == 4'h2;
  assign T41 = io_wb_req_ready & io_wb_req_valid;
  assign T42 = T63 & T43;
  assign T43 = T52 ? T49 : T44;
  assign T44 = T46 | T45;
  assign T45 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T46 = T48 | T47;
  assign T47 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T48 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T49 = T51 | T50;
  assign T50 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T51 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T52 = T54 | T53;
  assign T53 = io_req_bits_cmd == 5'h6;
  assign T54 = T56 | T55;
  assign T55 = io_req_bits_cmd == 5'h3;
  assign T56 = T60 | T57;
  assign T57 = T59 | T58;
  assign T58 = io_req_bits_cmd == 5'h4;
  assign T59 = io_req_bits_cmd[2'h3:2'h3];
  assign T60 = T62 | T61;
  assign T61 = io_req_bits_cmd == 5'h7;
  assign T62 = io_req_bits_cmd == 5'h1;
  assign T63 = T33 & io_req_bits_tag_match;
  assign T64 = T63 & T65;
  assign T65 = T43 ^ 1'h1;
  assign T66 = T67 ? 4'h1 : 4'h3;
  assign T67 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T68 = T33 & T69;
  assign T69 = io_req_bits_tag_match ^ 1'h1;
  assign T82 = T84 | T83;
  assign T83 = state == 4'h4;
  assign T84 = state == 4'h0;
  assign T205 = T207 & T206;
  assign T206 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T207 = wb_done | refill_done;
  assign wb_done = reply & T208;
  assign T208 = state == 4'h2;
  assign T209 = T86 ? 1'h0 : T210;
  assign T210 = T212 | T211;
  assign T211 = state == 4'h0;
  assign T212 = io_replay_ready & T213;
  assign T213 = state == 4'h8;
  assign T86 = io_meta_read_ready ^ 1'h1;
  assign T214 = T219 & T215;
  assign T215 = T216 ^ 1'h1;
  assign T216 = T218 | T217;
  assign T217 = io_req_bits_cmd == 5'h3;
  assign T218 = io_req_bits_cmd == 5'h2;
  assign T219 = T221 | T220;
  assign T220 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T156;
  assign T156 = T193 | T157;
  assign T157 = T190 & T158;
  assign T158 = T159 ^ 1'h1;
  assign T159 = T173 | T160;
  assign T160 = T162 & T161;
  assign T161 = io_mem_req_bits_a_type != 3'h1;
  assign T162 = T164 | T163;
  assign T163 = io_req_bits_cmd == 5'h6;
  assign T164 = T166 | T165;
  assign T165 = io_req_bits_cmd == 5'h3;
  assign T166 = T170 | T167;
  assign T167 = T169 | T168;
  assign T168 = io_req_bits_cmd == 5'h4;
  assign T169 = io_req_bits_cmd[2'h3:2'h3];
  assign T170 = T172 | T171;
  assign T171 = io_req_bits_cmd == 5'h7;
  assign T172 = io_req_bits_cmd == 5'h1;
  assign T173 = T183 & T174;
  assign T174 = T176 | T175;
  assign T175 = 3'h6 == io_mem_req_bits_a_type;
  assign T176 = T178 | T177;
  assign T177 = 3'h5 == io_mem_req_bits_a_type;
  assign T178 = T180 | T179;
  assign T179 = 3'h4 == io_mem_req_bits_a_type;
  assign T180 = T182 | T181;
  assign T181 = 3'h3 == io_mem_req_bits_a_type;
  assign T182 = 3'h2 == io_mem_req_bits_a_type;
  assign T183 = T187 | T184;
  assign T184 = T186 | T185;
  assign T185 = io_req_bits_cmd == 5'h4;
  assign T186 = io_req_bits_cmd[2'h3:2'h3];
  assign T187 = T189 | T188;
  assign T188 = io_req_bits_cmd == 5'h6;
  assign T189 = io_req_bits_cmd == 5'h0;
  assign T190 = T192 | T191;
  assign T191 = state == 4'h5;
  assign T192 = state == 4'h4;
  assign T193 = T195 | T194;
  assign T194 = state == 4'h3;
  assign T195 = T197 | T196;
  assign T196 = state == 4'h2;
  assign T197 = state == 4'h1;
  assign idx_match = req_idx == T74;
  assign T74 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T75 = T33 ? io_req_bits_addr : req_addr;
  assign T221 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T0;
  assign T0 = T73 | T1;
  assign T1 = T8 & T2;
  assign T2 = meta_hazard == 2'h0;
  assign T199 = reset ? 2'h0 : T3;
  assign T3 = T7 ? 2'h1 : T4;
  assign T4 = T6 ? T5 : meta_hazard;
  assign T5 = meta_hazard + 2'h1;
  assign T6 = meta_hazard != 2'h0;
  assign T7 = io_meta_write_ready & io_meta_write_valid;
  assign T8 = T70 & T9;
  assign T9 = state != 4'h3;
  assign T70 = T72 & T71;
  assign T71 = state != 4'h2;
  assign T72 = state != 4'h1;
  assign T73 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_master_xact_id = 3'h0;
  assign io_wb_req_bits_client_xact_id = 2'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T76 = T33 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = req_idx;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T77 = T33 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T78;
  assign T78 = T79 & ackq_io_enq_ready;
  assign T79 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T80;
  assign T80 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T85;
  assign T85 = T86 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_data = rpq_io_deq_bits_data;
  assign io_replay_bits_addr = T201;
  assign T201 = {12'h0, T87};
  assign T87 = T88;
  assign T88 = {io_tag, T89};
  assign T89 = {req_idx, T90};
  assign T90 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T91;
  assign T91 = T92 & rpq_io_deq_valid;
  assign T92 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T93;
  assign T93 = T113 ? meta_on_flush_state : line_state_state;
  assign T94 = T42 ? meta_on_hit_state : T95;
  assign T95 = T33 ? meta_on_flush_state : T96;
  assign T96 = T32 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T97;
  assign T97 = T104 ? 2'h1 : T98;
  assign T98 = T103 ? T101 : T99;
  assign T99 = T100 ? 2'h3 : 2'h0;
  assign T100 = io_mem_grant_bits_payload_g_type == 4'h5;
  assign T101 = T102 ? 2'h3 : 2'h2;
  assign T102 = io_mem_req_bits_a_type == 3'h1;
  assign T103 = io_mem_grant_bits_payload_g_type == 4'h2;
  assign T104 = io_mem_grant_bits_payload_g_type == 4'h1;
  assign meta_on_hit_state = T105;
  assign T105 = T106 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T106 = T110 | T107;
  assign T107 = T109 | T108;
  assign T108 = io_req_bits_cmd == 5'h4;
  assign T109 = io_req_bits_cmd[2'h3:2'h3];
  assign T110 = T112 | T111;
  assign T111 = io_req_bits_cmd == 5'h7;
  assign T112 = io_req_bits_cmd == 5'h1;
  assign meta_on_flush_state = 2'h0;
  assign T113 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T114;
  assign T114 = T116 | T115;
  assign T115 = state == 4'h3;
  assign T116 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T117;
  assign T117 = state == 4'h8;
  assign io_mem_resp_data = T202;
  assign T202 = {64'h0, req_data};
  assign T118 = T33 ? io_req_bits_data : req_data;
  assign io_mem_resp_addr = T119;
  assign T119 = T120 << 3'h4;
  assign T120 = {req_idx, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_a_type = acquire_type;
  assign T121 = T33 ? T136 : T122;
  assign T122 = T135 ? T123 : acquire_type;
  assign T123 = T124 ? 3'h1 : io_mem_req_bits_a_type;
  assign T124 = T126 | T125;
  assign T125 = io_req_bits_cmd == 5'h6;
  assign T126 = T128 | T127;
  assign T127 = io_req_bits_cmd == 5'h3;
  assign T128 = T132 | T129;
  assign T129 = T131 | T130;
  assign T130 = io_req_bits_cmd == 5'h4;
  assign T131 = io_req_bits_cmd[2'h3:2'h3];
  assign T132 = T134 | T133;
  assign T133 = io_req_bits_cmd == 5'h7;
  assign T134 = io_req_bits_cmd == 5'h1;
  assign T135 = io_req_sec_val & io_req_sec_rdy;
  assign T136 = T137 ? 3'h1 : 3'h0;
  assign T137 = T139 | T138;
  assign T138 = io_req_bits_cmd == 5'h6;
  assign T139 = T141 | T140;
  assign T140 = io_req_bits_cmd == 5'h3;
  assign T141 = T145 | T142;
  assign T142 = T144 | T143;
  assign T143 = io_req_bits_cmd == 5'h4;
  assign T144 = io_req_bits_cmd[2'h3:2'h3];
  assign T145 = T147 | T146;
  assign T146 = io_req_bits_cmd == 5'h7;
  assign T147 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_client_xact_id = 2'h1;
  assign io_mem_req_bits_addr = T148;
  assign T148 = T149;
  assign T149 = {io_tag, req_idx};
  assign io_mem_req_valid = T150;
  assign T150 = T151 & ackq_io_enq_ready;
  assign T151 = state == 4'h4;
  assign io_tag = T203;
  assign T203 = T152[5'h13:1'h0];
  assign T152 = req_addr >> 4'hc;
  assign io_idx_match = T153;
  assign T153 = T154 & idx_match;
  assign T154 = state != 4'h0;
  assign io_req_sec_rdy = T155;
  assign T155 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T198;
  assign T198 = state == 4'h0;
  Queue_14 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T214 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_data( io_req_bits_data ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_sdq_id ),
       .io_deq_ready( T209 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_data( rpq_io_deq_bits_data ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_11 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T205 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T204 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T68) begin
      state <= T66;
    end else if(T64) begin
      state <= 4'h4;
    end else if(T42) begin
      state <= 4'h6;
    end else if(T41) begin
      state <= 4'h2;
    end else if(T39) begin
      state <= 4'h3;
    end else if(T37) begin
      state <= 4'h4;
    end else if(T36) begin
      state <= 4'h5;
    end else if(T27) begin
      state <= 4'h6;
    end else if(T25) begin
      state <= 4'h7;
    end else if(T24) begin
      state <= 4'h8;
    end else if(T21) begin
      state <= 4'h0;
    end
    if(T33) begin
      refill_count <= 2'h0;
    end else if(T32) begin
      refill_count <= T31;
    end
    if(T33) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T7) begin
      meta_hazard <= 2'h1;
    end else if(T6) begin
      meta_hazard <= T5;
    end
    if(T33) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T33) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T42) begin
      line_state_state <= meta_on_hit_state;
    end else if(T33) begin
      line_state_state <= meta_on_flush_state;
    end else if(T32) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T33) begin
      req_data <= io_req_bits_data;
    end
    if(T33) begin
      acquire_type <= T136;
    end else if(T135) begin
      acquire_type <= T123;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[511:0] io_mem_req_bits_data,
    output[2:0] io_mem_req_bits_a_type,
    output[5:0] io_mem_req_bits_write_mask,
    output[2:0] io_mem_req_bits_subword_addr,
    output[3:0] io_mem_req_bits_atomic_opcode,
    output io_mem_resp_way_en,
    output[11:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire[4:0] T92;
  wire[4:0] T93;
  wire[4:0] T94;
  wire[4:0] T95;
  wire[4:0] T96;
  wire[4:0] T97;
  wire[4:0] T98;
  wire[4:0] T99;
  wire[4:0] T100;
  wire[4:0] T101;
  wire[4:0] T102;
  wire[4:0] T103;
  wire[4:0] T104;
  wire[4:0] T105;
  wire[4:0] T106;
  wire[4:0] T107;
  wire T108;
  wire[16:0] T21;
  wire[16:0] T22;
  reg [16:0] sdq_val;
  wire[16:0] T109;
  wire[31:0] T110;
  wire[31:0] T23;
  wire[31:0] T111;
  wire[31:0] T24;
  wire[31:0] T112;
  wire[16:0] T25;
  wire[16:0] T26;
  wire[16:0] T113;
  wire sdq_enq;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[16:0] T27;
  wire[16:0] T28;
  wire[16:0] T29;
  wire[16:0] T30;
  wire[16:0] T31;
  wire[16:0] T32;
  wire[16:0] T33;
  wire[16:0] T34;
  wire[16:0] T35;
  wire[16:0] T36;
  wire[16:0] T37;
  wire[16:0] T38;
  wire[16:0] T39;
  wire[16:0] T40;
  wire[16:0] T41;
  wire[16:0] T42;
  wire[16:0] T43;
  wire T44;
  wire[16:0] T45;
  wire[16:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire[31:0] T65;
  wire[31:0] T114;
  wire[16:0] T66;
  wire[16:0] T115;
  wire free_sdq;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[31:0] T75;
  wire[31:0] T116;
  wire T76;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T134;
  wire tag_match;
  wire[31:0] T88;
  wire[31:0] T133;
  wire[19:0] T89;
  wire[19:0] T90;
  wire[19:0] tagList_1;
  wire idxMatch_1;
  wire[19:0] T91;
  wire[19:0] tagList_0;
  wire idxMatch_0;
  wire T135;
  wire sdq_rdy;
  wire T85;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire idx_match;
  wire T140;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[63:0] T8;
  reg [63:0] sdq [16:0];
  wire[63:0] T9;
  wire T10;
  wire T11;
  wire[4:0] T12;
  reg [4:0] R77;
  wire[4:0] T78;
  wire[127:0] T79;
  wire[127:0] memRespMux_0_data;
  wire[127:0] memRespMux_1_data;
  wire T80;
  wire T132;
  wire[1:0] T81;
  wire[1:0] memRespMux_0_wmask;
  wire[1:0] memRespMux_1_wmask;
  wire[11:0] T82;
  wire[11:0] memRespMux_0_addr;
  wire[11:0] memRespMux_1_addr;
  wire T83;
  wire memRespMux_0_way_en;
  wire memRespMux_1_way_en;
  wire T84;
  wire T86;
  wire pri_rdy;
  wire T87;
  wire sec_rdy;
  wire meta_read_arb_io_in_1_ready;
  wire meta_read_arb_io_in_0_ready;
  wire meta_read_arb_io_out_valid;
  wire[5:0] meta_read_arb_io_out_bits_idx;
  wire[19:0] meta_read_arb_io_out_bits_tag;
  wire meta_write_arb_io_in_1_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_write_arb_io_out_valid;
  wire[5:0] meta_write_arb_io_out_bits_idx;
  wire meta_write_arb_io_out_bits_way_en;
  wire[19:0] meta_write_arb_io_out_bits_data_tag;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire mem_req_arb_io_in_1_ready;
  wire mem_req_arb_io_in_0_ready;
  wire mem_req_arb_io_out_valid;
  wire[25:0] mem_req_arb_io_out_bits_addr;
  wire[1:0] mem_req_arb_io_out_bits_client_xact_id;
  wire[511:0] mem_req_arb_io_out_bits_data;
  wire[2:0] mem_req_arb_io_out_bits_a_type;
  wire[5:0] mem_req_arb_io_out_bits_write_mask;
  wire[2:0] mem_req_arb_io_out_bits_subword_addr;
  wire[3:0] mem_req_arb_io_out_bits_atomic_opcode;
  wire mem_finish_arb_io_in_1_ready;
  wire mem_finish_arb_io_in_0_ready;
  wire mem_finish_arb_io_out_valid;
  wire[1:0] mem_finish_arb_io_out_bits_header_src;
  wire[1:0] mem_finish_arb_io_out_bits_header_dst;
  wire[2:0] mem_finish_arb_io_out_bits_payload_master_xact_id;
  wire wb_req_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire wb_req_arb_io_out_valid;
  wire[19:0] wb_req_arb_io_out_bits_tag;
  wire[5:0] wb_req_arb_io_out_bits_idx;
  wire wb_req_arb_io_out_bits_way_en;
  wire[1:0] wb_req_arb_io_out_bits_client_xact_id;
  wire[2:0] wb_req_arb_io_out_bits_master_xact_id;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire replay_arb_io_in_1_ready;
  wire replay_arb_io_in_0_ready;
  wire replay_arb_io_out_valid;
  wire replay_arb_io_out_bits_kill;
  wire[2:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_phys;
  wire[43:0] replay_arb_io_out_bits_addr;
  wire[7:0] replay_arb_io_out_bits_tag;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire MSHR_0_io_req_pri_rdy;
  wire MSHR_0_io_req_sec_rdy;
  wire MSHR_0_io_idx_match;
  wire[19:0] MSHR_0_io_tag;
  wire MSHR_0_io_mem_req_valid;
  wire[25:0] MSHR_0_io_mem_req_bits_addr;
  wire[1:0] MSHR_0_io_mem_req_bits_client_xact_id;
  wire[2:0] MSHR_0_io_mem_req_bits_a_type;
  wire MSHR_0_io_mem_resp_way_en;
  wire[11:0] MSHR_0_io_mem_resp_addr;
  wire[1:0] MSHR_0_io_mem_resp_wmask;
  wire[127:0] MSHR_0_io_mem_resp_data;
  wire MSHR_0_io_meta_read_valid;
  wire[5:0] MSHR_0_io_meta_read_bits_idx;
  wire[19:0] MSHR_0_io_meta_read_bits_tag;
  wire MSHR_0_io_meta_write_valid;
  wire[5:0] MSHR_0_io_meta_write_bits_idx;
  wire MSHR_0_io_meta_write_bits_way_en;
  wire[19:0] MSHR_0_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_0_io_meta_write_bits_data_coh_state;
  wire MSHR_0_io_replay_valid;
  wire MSHR_0_io_replay_bits_kill;
  wire[2:0] MSHR_0_io_replay_bits_typ;
  wire MSHR_0_io_replay_bits_phys;
  wire[43:0] MSHR_0_io_replay_bits_addr;
  wire[63:0] MSHR_0_io_replay_bits_data;
  wire[7:0] MSHR_0_io_replay_bits_tag;
  wire[4:0] MSHR_0_io_replay_bits_cmd;
  wire[4:0] MSHR_0_io_replay_bits_sdq_id;
  wire MSHR_0_io_mem_finish_valid;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_src;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_dst;
  wire[2:0] MSHR_0_io_mem_finish_bits_payload_master_xact_id;
  wire MSHR_0_io_wb_req_valid;
  wire[19:0] MSHR_0_io_wb_req_bits_tag;
  wire[5:0] MSHR_0_io_wb_req_bits_idx;
  wire MSHR_0_io_wb_req_bits_way_en;
  wire[1:0] MSHR_0_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_0_io_wb_req_bits_master_xact_id;
  wire[2:0] MSHR_0_io_wb_req_bits_r_type;
  wire MSHR_0_io_probe_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire MSHR_1_io_req_sec_rdy;
  wire MSHR_1_io_idx_match;
  wire[19:0] MSHR_1_io_tag;
  wire MSHR_1_io_mem_req_valid;
  wire[25:0] MSHR_1_io_mem_req_bits_addr;
  wire[1:0] MSHR_1_io_mem_req_bits_client_xact_id;
  wire[2:0] MSHR_1_io_mem_req_bits_a_type;
  wire MSHR_1_io_mem_resp_way_en;
  wire[11:0] MSHR_1_io_mem_resp_addr;
  wire[1:0] MSHR_1_io_mem_resp_wmask;
  wire[127:0] MSHR_1_io_mem_resp_data;
  wire MSHR_1_io_meta_read_valid;
  wire[5:0] MSHR_1_io_meta_read_bits_idx;
  wire[19:0] MSHR_1_io_meta_read_bits_tag;
  wire MSHR_1_io_meta_write_valid;
  wire[5:0] MSHR_1_io_meta_write_bits_idx;
  wire MSHR_1_io_meta_write_bits_way_en;
  wire[19:0] MSHR_1_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire MSHR_1_io_replay_valid;
  wire MSHR_1_io_replay_bits_kill;
  wire[2:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_phys;
  wire[43:0] MSHR_1_io_replay_bits_addr;
  wire[63:0] MSHR_1_io_replay_bits_data;
  wire[7:0] MSHR_1_io_replay_bits_tag;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire MSHR_1_io_mem_finish_valid;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_src;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_dst;
  wire[2:0] MSHR_1_io_mem_finish_bits_payload_master_xact_id;
  wire MSHR_1_io_wb_req_valid;
  wire[19:0] MSHR_1_io_wb_req_bits_tag;
  wire[5:0] MSHR_1_io_wb_req_bits_idx;
  wire MSHR_1_io_wb_req_bits_way_en;
  wire[1:0] MSHR_1_io_wb_req_bits_client_xact_id;
  wire[2:0] MSHR_1_io_wb_req_bits_master_xact_id;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire MSHR_1_io_probe_rdy;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R77 = {1{$random}};
  end
`endif

  assign T92 = T131 ? 1'h0 : T93;
  assign T93 = T130 ? 1'h1 : T94;
  assign T94 = T129 ? 2'h2 : T95;
  assign T95 = T128 ? 2'h3 : T96;
  assign T96 = T127 ? 3'h4 : T97;
  assign T97 = T126 ? 3'h5 : T98;
  assign T98 = T125 ? 3'h6 : T99;
  assign T99 = T124 ? 3'h7 : T100;
  assign T100 = T123 ? 4'h8 : T101;
  assign T101 = T122 ? 4'h9 : T102;
  assign T102 = T121 ? 4'ha : T103;
  assign T103 = T120 ? 4'hb : T104;
  assign T104 = T119 ? 4'hc : T105;
  assign T105 = T118 ? 4'hd : T106;
  assign T106 = T117 ? 4'he : T107;
  assign T107 = T108 ? 4'hf : 5'h10;
  assign T108 = T21[4'hf:4'hf];
  assign T21 = ~ T22;
  assign T22 = sdq_val[5'h10:1'h0];
  assign T109 = T110[5'h10:1'h0];
  assign T110 = reset ? 32'h0 : T23;
  assign T23 = T76 ? T24 : T111;
  assign T111 = {15'h0, sdq_val};
  assign T24 = T63 | T112;
  assign T112 = {15'h0, T25};
  assign T25 = T27 & T26;
  assign T26 = 17'h0 - T113;
  assign T113 = {16'h0, sdq_enq};
  assign sdq_enq = T20 & T13;
  assign T13 = T17 | T14;
  assign T14 = T16 | T15;
  assign T15 = io_req_bits_cmd == 5'h4;
  assign T16 = io_req_bits_cmd[2'h3:2'h3];
  assign T17 = T19 | T18;
  assign T18 = io_req_bits_cmd == 5'h7;
  assign T19 = io_req_bits_cmd == 5'h1;
  assign T20 = io_req_valid & io_req_ready;
  assign T27 = T62 ? 17'h1 : T28;
  assign T28 = T61 ? 17'h2 : T29;
  assign T29 = T60 ? 17'h4 : T30;
  assign T30 = T59 ? 17'h8 : T31;
  assign T31 = T58 ? 17'h10 : T32;
  assign T32 = T57 ? 17'h20 : T33;
  assign T33 = T56 ? 17'h40 : T34;
  assign T34 = T55 ? 17'h80 : T35;
  assign T35 = T54 ? 17'h100 : T36;
  assign T36 = T53 ? 17'h200 : T37;
  assign T37 = T52 ? 17'h400 : T38;
  assign T38 = T51 ? 17'h800 : T39;
  assign T39 = T50 ? 17'h1000 : T40;
  assign T40 = T49 ? 17'h2000 : T41;
  assign T41 = T48 ? 17'h4000 : T42;
  assign T42 = T47 ? 17'h8000 : T43;
  assign T43 = T44 ? 17'h10000 : 17'h0;
  assign T44 = T45[5'h10:5'h10];
  assign T45 = ~ T46;
  assign T46 = sdq_val[5'h10:1'h0];
  assign T47 = T45[4'hf:4'hf];
  assign T48 = T45[4'he:4'he];
  assign T49 = T45[4'hd:4'hd];
  assign T50 = T45[4'hc:4'hc];
  assign T51 = T45[4'hb:4'hb];
  assign T52 = T45[4'ha:4'ha];
  assign T53 = T45[4'h9:4'h9];
  assign T54 = T45[4'h8:4'h8];
  assign T55 = T45[3'h7:3'h7];
  assign T56 = T45[3'h6:3'h6];
  assign T57 = T45[3'h5:3'h5];
  assign T58 = T45[3'h4:3'h4];
  assign T59 = T45[2'h3:2'h3];
  assign T60 = T45[2'h2:2'h2];
  assign T61 = T45[1'h1:1'h1];
  assign T62 = T45[1'h0:1'h0];
  assign T63 = T116 & T64;
  assign T64 = ~ T65;
  assign T65 = T75 & T114;
  assign T114 = {15'h0, T66};
  assign T66 = 17'h0 - T115;
  assign T115 = {16'h0, free_sdq};
  assign free_sdq = T74 & T67;
  assign T67 = T71 | T68;
  assign T68 = T70 | T69;
  assign T69 = io_replay_bits_cmd == 5'h4;
  assign T70 = io_replay_bits_cmd[2'h3:2'h3];
  assign T71 = T73 | T72;
  assign T72 = io_replay_bits_cmd == 5'h7;
  assign T73 = io_replay_bits_cmd == 5'h1;
  assign T74 = io_replay_ready & io_replay_valid;
  assign T75 = 1'h1 << io_replay_bits_sdq_id;
  assign T116 = {15'h0, sdq_val};
  assign T76 = io_replay_valid | sdq_enq;
  assign T117 = T21[4'he:4'he];
  assign T118 = T21[4'hd:4'hd];
  assign T119 = T21[4'hc:4'hc];
  assign T120 = T21[4'hb:4'hb];
  assign T121 = T21[4'ha:4'ha];
  assign T122 = T21[4'h9:4'h9];
  assign T123 = T21[4'h8:4'h8];
  assign T124 = T21[3'h7:3'h7];
  assign T125 = T21[3'h6:3'h6];
  assign T126 = T21[3'h5:3'h5];
  assign T127 = T21[3'h4:3'h4];
  assign T128 = T21[2'h3:2'h3];
  assign T129 = T21[2'h2:2'h2];
  assign T130 = T21[1'h1:1'h1];
  assign T131 = T21[1'h0:1'h0];
  assign T134 = T135 & tag_match;
  assign tag_match = T133 == T88;
  assign T88 = io_req_bits_addr >> 4'hc;
  assign T133 = {12'h0, T89};
  assign T89 = T91 | T90;
  assign T90 = idxMatch_1 ? tagList_1 : 20'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T91 = idxMatch_0 ? tagList_0 : 20'h0;
  assign tagList_0 = MSHR_0_io_tag;
  assign idxMatch_0 = MSHR_0_io_idx_match;
  assign T135 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T85 ^ 1'h1;
  assign T85 = sdq_val == 17'h1ffff;
  assign T136 = T137 & tag_match;
  assign T137 = io_req_valid & sdq_rdy;
  assign T138 = T140 & T139;
  assign T139 = idx_match ^ 1'h1;
  assign idx_match = MSHR_0_io_idx_match | MSHR_1_io_idx_match;
  assign T140 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T0;
  assign T0 = T3 ? 1'h0 : T1;
  assign T1 = T2 == 1'h0;
  assign T2 = MSHR_0_io_req_pri_rdy ^ 1'h1;
  assign T3 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign io_probe_rdy = T4;
  assign T4 = T7 ? 1'h0 : T5;
  assign T5 = T6 == 1'h0;
  assign T6 = MSHR_0_io_probe_rdy ^ 1'h1;
  assign T7 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_master_xact_id = wb_req_arb_io_out_bits_master_xact_id;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_idx = wb_req_arb_io_out_bits_idx;
  assign io_wb_req_bits_tag = wb_req_arb_io_out_bits_tag;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_mem_finish_bits_payload_master_xact_id = mem_finish_arb_io_out_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mem_finish_arb_io_out_bits_header_dst;
  assign io_mem_finish_bits_header_src = mem_finish_arb_io_out_bits_header_src;
  assign io_mem_finish_valid = mem_finish_arb_io_out_valid;
  assign io_replay_bits_sdq_id = replay_arb_io_out_bits_sdq_id;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_data = T8;
  assign T8 = sdq[R77];
  assign T10 = sdq_enq & T11;
  assign T11 = T12 < 5'h11;
  assign T12 = T92[3'h4:1'h0];
  assign T78 = free_sdq ? replay_arb_io_out_bits_sdq_id : R77;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_mem_resp_data = T79;
  assign T79 = T80 ? memRespMux_1_data : memRespMux_0_data;
  assign memRespMux_0_data = MSHR_0_io_mem_resp_data;
  assign memRespMux_1_data = MSHR_1_io_mem_resp_data;
  assign T80 = T132;
  assign T132 = io_mem_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_mem_resp_wmask = T81;
  assign T81 = T80 ? memRespMux_1_wmask : memRespMux_0_wmask;
  assign memRespMux_0_wmask = MSHR_0_io_mem_resp_wmask;
  assign memRespMux_1_wmask = MSHR_1_io_mem_resp_wmask;
  assign io_mem_resp_addr = T82;
  assign T82 = T80 ? memRespMux_1_addr : memRespMux_0_addr;
  assign memRespMux_0_addr = MSHR_0_io_mem_resp_addr;
  assign memRespMux_1_addr = MSHR_1_io_mem_resp_addr;
  assign io_mem_resp_way_en = T83;
  assign T83 = T80 ? memRespMux_1_way_en : memRespMux_0_way_en;
  assign memRespMux_0_way_en = MSHR_0_io_mem_resp_way_en;
  assign memRespMux_1_way_en = MSHR_1_io_mem_resp_way_en;
  assign io_mem_req_bits_atomic_opcode = mem_req_arb_io_out_bits_atomic_opcode;
  assign io_mem_req_bits_subword_addr = mem_req_arb_io_out_bits_subword_addr;
  assign io_mem_req_bits_write_mask = mem_req_arb_io_out_bits_write_mask;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr = mem_req_arb_io_out_bits_addr;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign io_req_ready = T84;
  assign T84 = T86 & sdq_rdy;
  assign T86 = idx_match ? T87 : pri_rdy;
  assign pri_rdy = MSHR_0_io_req_pri_rdy | MSHR_1_io_req_pri_rdy;
  assign T87 = tag_match & sec_rdy;
  assign sec_rdy = MSHR_0_io_req_sec_rdy | MSHR_1_io_req_sec_rdy;
  Arbiter_6 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_in_0_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  Arbiter_7 mem_req_arb(
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       //.io_in_1_bits_data(  )
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       //.io_in_1_bits_write_mask(  )
       //.io_in_1_bits_subword_addr(  )
       //.io_in_1_bits_atomic_opcode(  )
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_req_valid ),
       .io_in_0_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       //.io_in_0_bits_data(  )
       .io_in_0_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       //.io_in_0_bits_write_mask(  )
       //.io_in_0_bits_subword_addr(  )
       //.io_in_0_bits_atomic_opcode(  )
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr( mem_req_arb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_write_mask( mem_req_arb_io_out_bits_write_mask ),
       .io_out_bits_subword_addr( mem_req_arb_io_out_bits_subword_addr ),
       .io_out_bits_atomic_opcode( mem_req_arb_io_out_bits_atomic_opcode )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign mem_req_arb.io_in_1_bits_data = {16{$random}};
    assign mem_req_arb.io_in_1_bits_write_mask = {1{$random}};
    assign mem_req_arb.io_in_1_bits_subword_addr = {1{$random}};
    assign mem_req_arb.io_in_1_bits_atomic_opcode = {1{$random}};
    assign mem_req_arb.io_in_0_bits_data = {16{$random}};
    assign mem_req_arb.io_in_0_bits_write_mask = {1{$random}};
    assign mem_req_arb.io_in_0_bits_subword_addr = {1{$random}};
    assign mem_req_arb.io_in_0_bits_atomic_opcode = {1{$random}};
  `endif
  Arbiter_8 mem_finish_arb(
       .io_in_1_ready( mem_finish_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_finish_valid ),
       .io_in_1_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_in_1_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( mem_finish_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_finish_valid ),
       .io_in_0_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_in_0_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_mem_finish_ready ),
       .io_out_valid( mem_finish_arb_io_out_valid ),
       .io_out_bits_header_src( mem_finish_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( mem_finish_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( mem_finish_arb_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  Arbiter_5 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( MSHR_1_io_wb_req_bits_master_xact_id ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_wb_req_valid ),
       .io_in_0_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( MSHR_0_io_wb_req_bits_master_xact_id ),
       .io_in_0_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_tag( wb_req_arb_io_out_bits_tag ),
       .io_out_bits_idx( wb_req_arb_io_out_bits_idx ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( wb_req_arb_io_out_bits_master_xact_id ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  Arbiter_9 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_data( MSHR_1_io_replay_bits_data ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_replay_valid ),
       .io_in_0_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_in_0_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_in_0_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_in_0_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_in_0_bits_data( MSHR_0_io_replay_bits_data ),
       .io_in_0_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_in_0_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       //.io_out_bits_data(  )
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_10 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( T138 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  MSHR_0 MSHR_0(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_0_io_req_pri_rdy ),
       .io_req_sec_val( T136 ),
       .io_req_sec_rdy( MSHR_0_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_data( io_req_bits_data ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_sdq_id( T92 ),
       .io_idx_match( MSHR_0_io_idx_match ),
       .io_tag( MSHR_0_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_0_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       //.io_mem_req_bits_data(  )
       .io_mem_req_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       //.io_mem_req_bits_write_mask(  )
       //.io_mem_req_bits_subword_addr(  )
       //.io_mem_req_bits_atomic_opcode(  )
       .io_mem_resp_way_en( MSHR_0_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_0_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_0_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_0_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_0_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_0_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_0_io_replay_valid ),
       .io_replay_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_replay_bits_data( MSHR_0_io_replay_bits_data ),
       .io_replay_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_0_ready ),
       .io_mem_finish_valid( MSHR_0_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_0_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( MSHR_0_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_0_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_0.io_mem_resp_wmask = {1{$random}};
  `endif
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T134 ),
       .io_req_sec_rdy( MSHR_1_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_data( io_req_bits_data ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_sdq_id( T92 ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       //.io_mem_req_bits_data(  )
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       //.io_mem_req_bits_write_mask(  )
       //.io_mem_req_bits_subword_addr(  )
       //.io_mem_req_bits_atomic_opcode(  )
       .io_mem_resp_way_en( MSHR_1_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_1_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_1_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_1_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_data( MSHR_1_io_replay_bits_data ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_1_ready ),
       .io_mem_finish_valid( MSHR_1_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( MSHR_1_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_1.io_mem_resp_wmask = {1{$random}};
  `endif

  always @(posedge clk) begin
    sdq_val <= T109;
    if (T10)
      sdq[T92] <= io_req_bits_data;
    if(free_sdq) begin
      R77 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [5:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [5:0] io_write_bits_idx,
    input  io_write_bits_way_en,
    input [19:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[19:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state
);

  wire[1:0] T0;
  wire[21:0] T1;
  wire[21:0] tags;
  wire[21:0] T2;
  wire[21:0] T3;
  wire[21:0] T4;
  wire[21:0] T20;
  wire T5;
  wire wmask;
  wire rst;
  reg [6:0] rst_cnt;
  wire[6:0] T21;
  wire[6:0] T6;
  wire[6:0] T7;
  wire[21:0] wdata;
  wire[21:0] T8;
  wire[1:0] T9;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T10;
  wire[19:0] T11;
  wire[19:0] rstVal_tag;
  wire T12;
  wire[5:0] T22;
  wire[6:0] waddr;
  wire[6:0] T23;
  reg [5:0] R13;
  wire[5:0] T14;
  wire[19:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    rst_cnt = {1{$random}};
    R13 = {1{$random}};
  end
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = tags[5'h15:1'h0];
  MetadataArray_tag_arr tag_arr (
    .CLK(clk),
    .W0A(T22),
    .W0E(T12),
    .W0I(wdata),
    .W0M(T3),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(tags)
  );
  assign T3 = T4;
  assign T4 = 22'h0 - T20;
  assign T20 = {21'h0, T5};
  assign T5 = wmask;
  assign wmask = rst ? 1'h1 : io_write_bits_way_en;
  assign rst = rst_cnt < 7'h40;
  assign T21 = reset ? 7'h0 : T6;
  assign T6 = rst ? T7 : rst_cnt;
  assign T7 = rst_cnt + 7'h1;
  assign wdata = T8;
  assign T8 = {T11, T9};
  assign T9 = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign rstVal_coh_state = T10;
  assign T10 = 2'h0;
  assign T11 = rst ? rstVal_tag : io_write_bits_data_tag;
  assign rstVal_tag = 20'h0;
  assign T12 = rst | io_write_valid;
  assign T22 = waddr[3'h5:1'h0];
  assign waddr = rst ? rst_cnt : T23;
  assign T23 = {1'h0, io_write_bits_idx};
  assign T14 = io_read_valid ? io_read_bits_idx : R13;
  assign io_resp_0_tag = T15;
  assign T15 = T1[5'h15:2'h2];
  assign io_write_ready = T16;
  assign T16 = rst ^ 1'h1;
  assign io_read_ready = T17;
  assign T17 = T19 & T18;
  assign T18 = io_write_valid ^ 1'h1;
  assign T19 = rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else if(rst) begin
      rst_cnt <= T7;
    end
    if(io_read_valid) begin
      R13 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_0(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [5:0] io_in_4_bits_idx,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [5:0] io_in_3_bits_idx,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [5:0] io_in_2_bits_idx,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[5:0] T5;
  wire[5:0] T6;
  wire[5:0] T7;
  wire T8;
  wire[2:0] T9;
  wire[5:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_idx = T5;
  assign T5 = T13 ? io_in_4_bits_idx : T6;
  assign T6 = T12 ? T10 : T7;
  assign T7 = T8 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T0;
  assign T10 = T11 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T11 = T9[1'h0:1'h0];
  assign T12 = T9[1'h1:1'h1];
  assign T13 = T9[2'h2:2'h2];
  assign io_out_valid = T14;
  assign T14 = T21 ? io_in_4_valid : T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T24;
  assign T24 = T25 & io_out_ready;
  assign T25 = T26 ^ 1'h1;
  assign T26 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T30 | io_in_2_valid;
  assign T30 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T34 | io_in_3_valid;
  assign T34 = T35 | io_in_2_valid;
  assign T35 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input  io_read_bits_way_en,
    input [11:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input  io_write_bits_way_en,
    input [11:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [127:0] io_write_bits_data,
    output[127:0] io_resp_0
);

  wire[127:0] T0;
  wire T12;
  wire[7:0] raddr;
  wire[127:0] T2;
  wire[127:0] T3;
  wire[127:0] T4;
  wire[63:0] T5;
  wire[63:0] T13;
  wire T6;
  wire[63:0] T7;
  wire[63:0] T14;
  wire T8;
  wire T9;
  wire[7:0] waddr;
  reg [7:0] R10;
  wire[7:0] T11;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R10 = {1{$random}};
  end
`endif

  assign io_resp_0 = T0;
  assign T12 = io_read_bits_way_en & io_read_valid;
  assign raddr = io_read_bits_addr >> 3'h4;
  DataArray_T1 T1 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T9),
    .W0I(io_write_bits_data),
    .W0M(T3),
    .R1A(raddr),
    .R1E(T12),
    .R1O(T0)
  );
  assign T3 = T4;
  assign T4 = {T7, T5};
  assign T5 = 64'h0 - T13;
  assign T13 = {63'h0, T6};
  assign T6 = io_write_bits_wmask[1'h0:1'h0];
  assign T7 = 64'h0 - T14;
  assign T14 = {63'h0, T8};
  assign T8 = io_write_bits_wmask[1'h1:1'h1];
  assign T9 = io_write_bits_way_en & io_write_valid;
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T11 = T12 ? raddr : R10;
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T12) begin
      R10 <= raddr;
    end
  end
endmodule

module Arbiter_2(
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits_way_en,
    input [11:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits_way_en,
    input [11:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[11:0] T4;
  wire[11:0] T5;
  wire T6;
  wire[1:0] T7;
  wire[11:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : T3;
  assign T3 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = T0;
  assign T8 = T9 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T9 = T7[1'h0:1'h0];
  assign T10 = T7[1'h1:1'h1];
  assign io_out_bits_way_en = T11;
  assign T11 = T16 ? T14 : T12;
  assign T12 = T13 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T13 = T7[1'h0:1'h0];
  assign T14 = T15 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T15 = T7[1'h0:1'h0];
  assign T16 = T7[1'h1:1'h1];
  assign io_out_valid = T17;
  assign T17 = T22 ? T20 : T18;
  assign T18 = T19 ? io_in_1_valid : io_in_0_valid;
  assign T19 = T7[1'h0:1'h0];
  assign T20 = T21 ? io_in_3_valid : io_in_2_valid;
  assign T21 = T7[1'h0:1'h0];
  assign T22 = T7[1'h1:1'h1];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T25;
  assign T25 = T26 & io_out_ready;
  assign T26 = T27 ^ 1'h1;
  assign T27 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 | io_in_2_valid;
  assign T31 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[127:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[11:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T2;
  assign T2 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T3 = T0;
  assign io_out_bits_wmask = T4;
  assign T4 = T3 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T5;
  assign T5 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T6;
  assign T6 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [3:0] io_cmd,
    input [2:0] io_typ,
    input [63:0] io_lhs,
    input [63:0] io_rhs,
    output[63:0] io_out
);

  wire[63:0] T118;
  wire[87:0] T0;
  wire[87:0] T1;
  wire[87:0] T119;
  wire[87:0] T2;
  wire[87:0] wmask;
  wire[87:0] T3;
  wire[47:0] T4;
  wire[23:0] T5;
  wire[15:0] T6;
  wire[7:0] T7;
  wire[7:0] T120;
  wire T8;
  wire[10:0] T9;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[10:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[10:0] T121;
  wire[8:0] T18;
  wire[2:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[10:0] T122;
  wire[7:0] T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T123;
  wire T30;
  wire[7:0] T31;
  wire[7:0] T124;
  wire T32;
  wire[23:0] T33;
  wire[15:0] T34;
  wire[7:0] T35;
  wire[7:0] T125;
  wire T36;
  wire[7:0] T37;
  wire[7:0] T126;
  wire T38;
  wire[7:0] T39;
  wire[7:0] T127;
  wire T40;
  wire[39:0] T41;
  wire[23:0] T42;
  wire[15:0] T43;
  wire[7:0] T44;
  wire[7:0] T128;
  wire T45;
  wire[7:0] T46;
  wire[7:0] T129;
  wire T47;
  wire[7:0] T48;
  wire[7:0] T130;
  wire T49;
  wire[15:0] T50;
  wire[7:0] T51;
  wire[7:0] T131;
  wire T52;
  wire[7:0] T53;
  wire[7:0] T132;
  wire T54;
  wire[87:0] T55;
  wire[87:0] T133;
  wire[63:0] out;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  wire[63:0] T60;
  wire[63:0] T61;
  wire[63:0] rhs;
  wire[63:0] T62;
  wire[31:0] T63;
  wire[63:0] T64;
  wire[31:0] T65;
  wire[15:0] T66;
  wire[63:0] T67;
  wire[31:0] T68;
  wire[15:0] T69;
  wire[7:0] T70;
  wire T71;
  wire max;
  wire T72;
  wire[4:0] T134;
  wire T73;
  wire[4:0] T135;
  wire min;
  wire T74;
  wire[4:0] T136;
  wire T75;
  wire[4:0] T137;
  wire less;
  wire T76;
  wire cmp_rhs;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire word;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire cmp_lhs;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire sgned;
  wire T93;
  wire[4:0] T138;
  wire T94;
  wire[4:0] T139;
  wire lt;
  wire T95;
  wire T96;
  wire lt_lo;
  wire[31:0] T97;
  wire[31:0] T98;
  wire eq_hi;
  wire[31:0] T99;
  wire[31:0] T100;
  wire lt_hi;
  wire[31:0] T101;
  wire[31:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire[63:0] T106;
  wire T107;
  wire[4:0] T140;
  wire[63:0] T108;
  wire T109;
  wire[4:0] T141;
  wire[63:0] T110;
  wire T111;
  wire[4:0] T142;
  wire[63:0] adder_out;
  wire[63:0] T112;
  wire[63:0] mask;
  wire[63:0] T143;
  wire[31:0] T113;
  wire T114;
  wire[63:0] T115;
  wire[63:0] T116;
  wire T117;
  wire[4:0] T144;


  assign io_out = T118;
  assign T118 = T0[6'h3f:1'h0];
  assign T0 = T55 | T1;
  assign T1 = T2 & T119;
  assign T119 = {24'h0, io_lhs};
  assign T2 = ~ wmask;
  assign wmask = T3;
  assign T3 = {T41, T4};
  assign T4 = {T33, T5};
  assign T5 = {T31, T6};
  assign T6 = {T29, T7};
  assign T7 = 8'h0 - T120;
  assign T120 = {7'h0, T8};
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T26 ? T122 : T10;
  assign T10 = T21 ? T121 : T11;
  assign T11 = T15 ? T12 : 11'hff;
  assign T12 = 4'hf << T13;
  assign T13 = {T14, 2'h0};
  assign T14 = io_addr[2'h2:2'h2];
  assign T15 = T17 | T16;
  assign T16 = io_typ == 3'h6;
  assign T17 = io_typ == 3'h2;
  assign T121 = {2'h0, T18};
  assign T18 = 2'h3 << T19;
  assign T19 = {T20, 1'h0};
  assign T20 = io_addr[2'h2:1'h1];
  assign T21 = T23 | T22;
  assign T22 = io_typ == 3'h5;
  assign T23 = io_typ == 3'h1;
  assign T122 = {3'h0, T24};
  assign T24 = 1'h1 << T25;
  assign T25 = io_addr[2'h2:1'h0];
  assign T26 = T28 | T27;
  assign T27 = io_typ == 3'h4;
  assign T28 = io_typ == 3'h0;
  assign T29 = 8'h0 - T123;
  assign T123 = {7'h0, T30};
  assign T30 = T9[1'h1:1'h1];
  assign T31 = 8'h0 - T124;
  assign T124 = {7'h0, T32};
  assign T32 = T9[2'h2:2'h2];
  assign T33 = {T39, T34};
  assign T34 = {T37, T35};
  assign T35 = 8'h0 - T125;
  assign T125 = {7'h0, T36};
  assign T36 = T9[2'h3:2'h3];
  assign T37 = 8'h0 - T126;
  assign T126 = {7'h0, T38};
  assign T38 = T9[3'h4:3'h4];
  assign T39 = 8'h0 - T127;
  assign T127 = {7'h0, T40};
  assign T40 = T9[3'h5:3'h5];
  assign T41 = {T50, T42};
  assign T42 = {T48, T43};
  assign T43 = {T46, T44};
  assign T44 = 8'h0 - T128;
  assign T128 = {7'h0, T45};
  assign T45 = T9[3'h6:3'h6];
  assign T46 = 8'h0 - T129;
  assign T129 = {7'h0, T47};
  assign T47 = T9[3'h7:3'h7];
  assign T48 = 8'h0 - T130;
  assign T130 = {7'h0, T49};
  assign T49 = T9[4'h8:4'h8];
  assign T50 = {T53, T51};
  assign T51 = 8'h0 - T131;
  assign T131 = {7'h0, T52};
  assign T52 = T9[4'h9:4'h9];
  assign T53 = 8'h0 - T132;
  assign T132 = {7'h0, T54};
  assign T54 = T9[4'ha:4'ha];
  assign T55 = wmask & T133;
  assign T133 = {24'h0, out};
  assign out = T117 ? adder_out : T56;
  assign T56 = T111 ? T110 : T57;
  assign T57 = T109 ? T108 : T58;
  assign T58 = T107 ? T106 : T59;
  assign T59 = T71 ? io_lhs : T60;
  assign T60 = T26 ? T67 : T61;
  assign T61 = T21 ? T64 : rhs;
  assign rhs = T15 ? T62 : io_rhs;
  assign T62 = {T63, T63};
  assign T63 = io_rhs[5'h1f:1'h0];
  assign T64 = {T65, T65};
  assign T65 = {T66, T66};
  assign T66 = io_rhs[4'hf:1'h0];
  assign T67 = {T68, T68};
  assign T68 = {T69, T69};
  assign T69 = {T70, T70};
  assign T70 = io_rhs[3'h7:1'h0];
  assign T71 = less ? min : max;
  assign max = T73 | T72;
  assign T72 = T134 == 5'hf;
  assign T134 = {1'h0, io_cmd};
  assign T73 = T135 == 5'hd;
  assign T135 = {1'h0, io_cmd};
  assign min = T75 | T74;
  assign T74 = T136 == 5'he;
  assign T136 = {1'h0, io_cmd};
  assign T75 = T137 == 5'hc;
  assign T137 = {1'h0, io_cmd};
  assign less = T105 ? lt : T76;
  assign T76 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T79 ? T78 : T77;
  assign T77 = rhs[6'h3f:6'h3f];
  assign T78 = rhs[5'h1f:5'h1f];
  assign T79 = word & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = io_addr[2'h2:2'h2];
  assign word = T83 | T82;
  assign T82 = io_typ == 3'h4;
  assign T83 = T85 | T84;
  assign T84 = io_typ == 3'h0;
  assign T85 = T87 | T86;
  assign T86 = io_typ == 3'h6;
  assign T87 = io_typ == 3'h2;
  assign cmp_lhs = T90 ? T89 : T88;
  assign T88 = io_lhs[6'h3f:6'h3f];
  assign T89 = io_lhs[5'h1f:5'h1f];
  assign T90 = word & T91;
  assign T91 = T92 ^ 1'h1;
  assign T92 = io_addr[2'h2:2'h2];
  assign sgned = T94 | T93;
  assign T93 = T138 == 5'hd;
  assign T138 = {1'h0, io_cmd};
  assign T94 = T139 == 5'hc;
  assign T139 = {1'h0, io_cmd};
  assign lt = word ? T103 : T95;
  assign T95 = lt_hi | T96;
  assign T96 = eq_hi & lt_lo;
  assign lt_lo = T98 < T97;
  assign T97 = rhs[5'h1f:1'h0];
  assign T98 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T100 == T99;
  assign T99 = rhs[6'h3f:6'h20];
  assign T100 = io_lhs[6'h3f:6'h20];
  assign lt_hi = T102 < T101;
  assign T101 = rhs[6'h3f:6'h20];
  assign T102 = io_lhs[6'h3f:6'h20];
  assign T103 = T104 ? lt_hi : lt_lo;
  assign T104 = io_addr[2'h2:2'h2];
  assign T105 = cmp_lhs == cmp_rhs;
  assign T106 = io_lhs ^ rhs;
  assign T107 = T140 == 5'h9;
  assign T140 = {1'h0, io_cmd};
  assign T108 = io_lhs | rhs;
  assign T109 = T141 == 5'ha;
  assign T141 = {1'h0, io_cmd};
  assign T110 = io_lhs & rhs;
  assign T111 = T142 == 5'hb;
  assign T142 = {1'h0, io_cmd};
  assign adder_out = T115 + T112;
  assign T112 = rhs & mask;
  assign mask = 64'hffffffffffffffff ^ T143;
  assign T143 = {32'h0, T113};
  assign T113 = T114 << 5'h1f;
  assign T114 = io_addr[2'h2:2'h2];
  assign T115 = T116;
  assign T116 = io_lhs & mask;
  assign T117 = T144 == 5'h8;
  assign T144 = {1'h0, io_cmd};
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_master_xact_id,
    input [511:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_master_xact_id,
    input [511:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_master_xact_id,
    output[511:0] io_out_bits_data,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[511:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire[25:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_data = T4;
  assign T4 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_master_xact_id = T5;
  assign T5 = T3 ? io_in_1_bits_master_xact_id : io_in_0_bits_master_xact_id;
  assign io_out_bits_client_xact_id = T6;
  assign T6 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T7;
  assign T7 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T8;
  assign T8 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module FlowThroughSerializer_0(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [1:0] io_in_bits_payload_client_xact_id,
    input [2:0] io_in_bits_payload_master_xact_id,
    input [3:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  active;
  wire T46;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T47;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire[1:0] T48;
  wire[1:0] T18;
  wire T19;
  wire[3:0] T20;
  reg [3:0] rbits_payload_g_type;
  wire[3:0] T49;
  wire[3:0] T21;
  wire[2:0] T22;
  reg [2:0] rbits_payload_master_xact_id;
  wire[2:0] T50;
  wire[2:0] T23;
  wire[1:0] T24;
  reg [1:0] rbits_payload_client_xact_id;
  wire[1:0] T51;
  wire[1:0] T25;
  wire[511:0] T26;
  wire[511:0] T27;
  reg [511:0] rbits_payload_data;
  wire[511:0] T52;
  wire[511:0] T28;
  wire[511:0] T53;
  wire[127:0] T29;
  wire[127:0] T30;
  wire[127:0] shifter_0;
  wire[127:0] T31;
  wire[127:0] shifter_1;
  wire[127:0] T32;
  wire T33;
  wire[1:0] T34;
  wire[127:0] T35;
  wire[127:0] shifter_2;
  wire[127:0] T36;
  wire[127:0] shifter_3;
  wire[127:0] T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  reg [1:0] rbits_header_dst;
  wire[1:0] T54;
  wire[1:0] T41;
  wire[1:0] T42;
  reg [1:0] rbits_header_src;
  wire[1:0] T55;
  wire[1:0] T43;
  wire T44;
  wire T45;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    active = {1{$random}};
    cnt = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T14 ? 1'h1 : T1;
  assign T1 = T6 ? T2 : 1'h0;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 | T4;
  assign T4 = io_in_bits_payload_g_type == 4'h2;
  assign T5 = io_in_bits_payload_g_type == 4'h1;
  assign T6 = T7 & io_in_valid;
  assign T7 = active ^ 1'h1;
  assign T46 = reset ? 1'h0 : T8;
  assign T8 = T14 ? 1'h0 : T9;
  assign T9 = T10 ? 1'h1 : active;
  assign T10 = T6 & T11;
  assign T11 = T13 | T12;
  assign T12 = io_in_bits_payload_g_type == 4'h2;
  assign T13 = io_in_bits_payload_g_type == 4'h1;
  assign T14 = T19 & wrap;
  assign wrap = cnt == 2'h3;
  assign T47 = reset ? 2'h0 : T15;
  assign T15 = T14 ? 2'h0 : T16;
  assign T16 = T19 ? T18 : T17;
  assign T17 = T10 ? T48 : cnt;
  assign T48 = {1'h0, io_out_ready};
  assign T18 = cnt + 2'h1;
  assign T19 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T20;
  assign T20 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T49 = reset ? io_in_bits_payload_g_type : T21;
  assign T21 = T10 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_master_xact_id = T22;
  assign T22 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T50 = reset ? io_in_bits_payload_master_xact_id : T23;
  assign T23 = T10 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T24;
  assign T24 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T51 = reset ? io_in_bits_payload_client_xact_id : T25;
  assign T25 = T10 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T26;
  assign T26 = active ? T53 : T27;
  assign T27 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T52 = reset ? io_in_bits_payload_data : T28;
  assign T28 = T10 ? io_in_bits_payload_data : rbits_payload_data;
  assign T53 = {384'h0, T29};
  assign T29 = T39 ? T35 : T30;
  assign T30 = T33 ? shifter_1 : shifter_0;
  assign shifter_0 = T31;
  assign T31 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T32;
  assign T32 = rbits_payload_data[8'hff:8'h80];
  assign T33 = T34[1'h0:1'h0];
  assign T34 = cnt;
  assign T35 = T38 ? shifter_3 : shifter_2;
  assign shifter_2 = T36;
  assign T36 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T37;
  assign T37 = rbits_payload_data[9'h1ff:9'h180];
  assign T38 = T34[1'h0:1'h0];
  assign T39 = T34[1'h1:1'h1];
  assign io_out_bits_header_dst = T40;
  assign T40 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T54 = reset ? io_in_bits_header_dst : T41;
  assign T41 = T10 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T42;
  assign T42 = active ? rbits_header_src : io_in_bits_header_src;
  assign T55 = reset ? io_in_bits_header_src : T43;
  assign T43 = T10 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T44;
  assign T44 = active | io_in_valid;
  assign io_in_ready = T45;
  assign T45 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      active <= 1'h0;
    end else if(T14) begin
      active <= 1'h0;
    end else if(T10) begin
      active <= 1'h1;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T14) begin
      cnt <= 2'h0;
    end else if(T19) begin
      cnt <= T18;
    end else if(T10) begin
      cnt <= T48;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T10) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T10) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T10) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T10) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T10) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T10) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input  io_cpu_req_bits_kill,
    input [2:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_phys,
    input [43:0] io_cpu_req_bits_addr,
    input [63:0] io_cpu_req_bits_data,
    input [7:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    output io_cpu_resp_valid,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output[2:0] io_cpu_resp_bits_typ,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data,
    output[63:0] io_cpu_resp_bits_data_subword,
    output[7:0] io_cpu_resp_bits_tag,
    output[3:0] io_cpu_resp_bits_cmd,
    output[43:0] io_cpu_resp_bits_addr,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[7:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    output io_cpu_ordered,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [2:0] io_mem_probe_bits_payload_master_xact_id,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[1:0] io_mem_release_bits_header_src,
    output[1:0] io_mem_release_bits_header_dst,
    output[25:0] io_mem_release_bits_payload_addr,
    output[1:0] io_mem_release_bits_payload_client_xact_id,
    output[2:0] io_mem_release_bits_payload_master_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type
);

  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  reg [63:0] s2_req_data;
  wire[63:0] T161;
  wire[63:0] T162;
  wire[63:0] T163;
  reg  s1_replay;
  wire T343;
  wire T26;
  wire T164;
  wire s1_write;
  wire T119;
  wire T120;
  reg [4:0] s1_req_cmd;
  wire[4:0] T19;
  wire[4:0] T20;
  wire[4:0] T21;
  reg [4:0] s2_req_cmd;
  wire[4:0] T18;
  wire s2_recycle;
  wire T22;
  reg  s2_recycle_next;
  wire T342;
  wire T23;
  wire T24;
  wire T25;
  reg  s1_valid;
  wire T344;
  wire T27;
  wire T28;
  wire s2_recycle_ecc;
  wire s2_data_correctable;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire s2_word_idx;
  reg [43:0] s2_req_addr;
  wire[43:0] T33;
  wire[43:0] T345;
  wire[31:0] s1_addr;
  wire[12:0] T34;
  reg [43:0] s1_req_addr;
  wire[43:0] T35;
  wire[43:0] T36;
  wire[43:0] T37;
  wire[43:0] T38;
  wire[43:0] T39;
  wire[43:0] T346;
  wire[31:0] T40;
  wire[25:0] T41;
  wire[43:0] T347;
  wire[31:0] T42;
  wire[25:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire s2_hit;
  wire T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  reg [1:0] s2_hit_state_state;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire s2_tag_match;
  reg  s2_tag_match_way;
  wire T79;
  wire s1_tag_match_way;
  wire T80;
  wire T81;
  wire T82;
  wire s1_tag_eq_way;
  wire T83;
  wire[19:0] T84;
  wire T85;
  wire s2_replay;
  wire T86;
  reg  R87;
  wire T348;
  reg  s2_valid;
  wire T349;
  wire s1_valid_masked;
  wire T88;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  reg  s1_clk_en;
  reg [63:0] s1_req_data;
  wire[63:0] T165;
  wire[63:0] T166;
  wire[63:0] T167;
  wire T168;
  reg  s1_recycled;
  wire T169;
  wire[63:0] T373;
  wire[127:0] s2_data_word;
  wire[127:0] s2_data_word_prebypass;
  wire[6:0] T186;
  wire[127:0] s2_data_uncorrected;
  wire[127:0] T187;
  wire[63:0] T188;
  wire[127:0] s2_data_0;
  wire[127:0] T189;
  wire[127:0] T190;
  reg [63:0] R191;
  wire[63:0] T352;
  wire[127:0] T192;
  wire[127:0] T353;
  wire[127:0] T193;
  wire T194;
  wire T195;
  reg [63:0] R196;
  wire[63:0] T197;
  wire[63:0] T198;
  wire[63:0] T199;
  wire[127:0] T354;
  reg [63:0] s2_store_bypass_data;
  wire[63:0] T200;
  wire[63:0] T201;
  wire[63:0] T202;
  reg [63:0] s4_req_data;
  wire[63:0] T203;
  wire T204;
  reg  s3_valid;
  wire T355;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire s2_sc_fail;
  wire T171;
  wire s2_lrsc_addr_match;
  wire T172;
  wire[37:0] T173;
  reg [37:0] lrsc_addr;
  wire[37:0] T174;
  wire[37:0] T175;
  wire T17;
  wire s2_lr;
  wire T89;
  wire T90;
  wire s2_valid_masked;
  wire T91;
  wire T92;
  wire s2_nack;
  wire s2_nack_miss;
  wire T93;
  wire T94;
  wire T95;
  wire s2_nack_victim;
  reg  s2_nack_hit;
  wire T96;
  wire s1_nack;
  wire T97;
  wire T98;
  wire T99;
  wire[5:0] T100;
  wire T101;
  wire T102;
  wire lrsc_valid;
  reg [4:0] lrsc_count;
  wire[4:0] T341;
  wire[4:0] T10;
  wire[4:0] T11;
  wire[4:0] T12;
  wire[4:0] T13;
  wire[4:0] T14;
  wire T15;
  wire T16;
  wire T103;
  wire s2_sc;
  wire T215;
  wire T216;
  reg [63:0] s3_req_data;
  wire[63:0] T356;
  wire[127:0] T217;
  wire[127:0] T357;
  wire[63:0] T218;
  wire[127:0] T219;
  wire[127:0] T358;
  wire[127:0] s2_data_corrected;
  wire[127:0] T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  reg [4:0] s3_req_cmd;
  wire[4:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire[40:0] T242;
  reg [43:0] s3_req_addr;
  wire[43:0] T243;
  wire[40:0] T359;
  wire[28:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire[40:0] T255;
  wire[40:0] T360;
  wire[28:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  reg [4:0] s4_req_cmd;
  wire[4:0] T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire[40:0] T273;
  reg [43:0] s4_req_addr;
  wire[43:0] T274;
  wire[40:0] T361;
  wire[28:0] T275;
  reg  s4_valid;
  wire T362;
  wire T276;
  reg  s2_store_bypass;
  wire T277;
  wire T278;
  reg [2:0] s2_req_typ;
  wire[2:0] T140;
  reg [2:0] s1_req_typ;
  wire[2:0] T137;
  wire[2:0] T138;
  wire[2:0] T139;
  wire[3:0] T374;
  wire[5:0] T375;
  wire[127:0] T376;
  wire[1:0] T377;
  wire T378;
  wire T379;
  wire[11:0] T380;
  reg  s3_way;
  wire T381;
  wire[127:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire[11:0] T389;
  wire[11:0] T390;
  wire[11:0] T391;
  wire[127:0] T392;
  wire[127:0] T393;
  wire[63:0] wdata_encoded_0;
  wire[63:0] wdata_encoded_1;
  wire[5:0] T394;
  wire[37:0] T395;
  wire[5:0] T396;
  wire[37:0] T397;
  reg  s1_req_phys;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  reg  s2_req_phys;
  wire T403;
  wire[30:0] T404;
  wire T405;
  wire T406;
  wire T407;
  wire s1_readwrite;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire s1_read;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T412;
  wire T413;
  wire T414;
  wire[1:0] T415;
  wire[1:0] s2_replaced_way_en;
  reg  R416;
  wire T417;
  wire[1:0] T418;
  wire[1:0] T419;
  reg [1:0] s2_repl_meta_coh_state;
  wire[1:0] T420;
  wire[1:0] T421;
  wire[19:0] T422;
  reg [19:0] s2_repl_meta_tag;
  wire[19:0] T423;
  wire[19:0] T424;
  reg [7:0] s2_req_tag;
  wire[7:0] T158;
  reg [7:0] s1_req_tag;
  wire[7:0] T155;
  wire[7:0] T156;
  wire[7:0] T157;
  reg  s2_req_kill;
  wire T425;
  reg  s1_req_kill;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[1:0] probe_bits_p_type;
  wire[2:0] probe_bits_master_xact_id;
  wire[25:0] probe_bits_addr;
  wire T452;
  wire T453;
  wire probe_valid;
  wire[2:0] T0;
  wire[511:0] T1;
  wire[2:0] T2;
  wire[1:0] T3;
  wire[25:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire probe_ready;
  wire T8;
  wire T9;
  wire[3:0] T104;
  wire[2:0] T105;
  wire[5:0] T106;
  wire[2:0] T107;
  wire[511:0] T108;
  wire[1:0] T109;
  wire[25:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T125;
  wire T132;
  wire misaligned;
  wire T133;
  wire T134;
  wire[2:0] T135;
  wire T136;
  wire T141;
  wire T142;
  wire T143;
  wire[1:0] T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T159;
  wire T160;
  wire s1_sc;
  wire[3:0] T350;
  wire[63:0] T170;
  wire[63:0] T351;
  wire[63:0] T176;
  wire[7:0] T177;
  wire[7:0] T178;
  wire[7:0] T179;
  wire[63:0] T180;
  wire[15:0] T181;
  wire[15:0] T182;
  wire[63:0] T183;
  wire[31:0] T184;
  wire[31:0] T185;
  wire[31:0] T279;
  wire T280;
  wire[31:0] T281;
  wire[31:0] T282;
  wire[31:0] T283;
  wire[31:0] T363;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire[15:0] T296;
  wire T297;
  wire[47:0] T298;
  wire[47:0] T299;
  wire[47:0] T300;
  wire[47:0] T364;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire[7:0] T306;
  wire T307;
  wire[55:0] T308;
  wire[55:0] T309;
  wire[55:0] T310;
  wire[55:0] T365;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  reg  block_miss;
  wire T366;
  wire T339;
  wire T340;
  wire wb_io_req_ready;
  wire wb_io_meta_read_valid;
  wire[5:0] wb_io_meta_read_bits_idx;
  wire[19:0] wb_io_meta_read_bits_tag;
  wire wb_io_data_req_valid;
  wire wb_io_data_req_bits_way_en;
  wire[11:0] wb_io_data_req_bits_addr;
  wire wb_io_release_valid;
  wire[25:0] wb_io_release_bits_addr;
  wire[1:0] wb_io_release_bits_client_xact_id;
  wire[2:0] wb_io_release_bits_master_xact_id;
  wire[511:0] wb_io_release_bits_data;
  wire[2:0] wb_io_release_bits_r_type;
  wire prober_io_req_ready;
  wire prober_io_rep_valid;
  wire[25:0] prober_io_rep_bits_addr;
  wire[1:0] prober_io_rep_bits_client_xact_id;
  wire[2:0] prober_io_rep_bits_master_xact_id;
  wire[511:0] prober_io_rep_bits_data;
  wire[2:0] prober_io_rep_bits_r_type;
  wire prober_io_meta_read_valid;
  wire[5:0] prober_io_meta_read_bits_idx;
  wire[19:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_write_valid;
  wire[5:0] prober_io_meta_write_bits_idx;
  wire prober_io_meta_write_bits_way_en;
  wire[19:0] prober_io_meta_write_bits_data_tag;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire prober_io_wb_req_valid;
  wire[19:0] prober_io_wb_req_bits_tag;
  wire[5:0] prober_io_wb_req_bits_idx;
  wire prober_io_wb_req_bits_way_en;
  wire[1:0] prober_io_wb_req_bits_client_xact_id;
  wire[2:0] prober_io_wb_req_bits_master_xact_id;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire meta_io_read_ready;
  wire meta_io_write_ready;
  wire[19:0] meta_io_resp_0_tag;
  wire[1:0] meta_io_resp_0_coh_state;
  wire metaReadArb_io_in_4_ready;
  wire metaReadArb_io_in_3_ready;
  wire metaReadArb_io_in_2_ready;
  wire metaReadArb_io_in_1_ready;
  wire metaReadArb_io_out_valid;
  wire[5:0] metaReadArb_io_out_bits_idx;
  wire metaWriteArb_io_in_1_ready;
  wire metaWriteArb_io_in_0_ready;
  wire metaWriteArb_io_out_valid;
  wire[5:0] metaWriteArb_io_out_bits_idx;
  wire metaWriteArb_io_out_bits_way_en;
  wire[19:0] metaWriteArb_io_out_bits_data_tag;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire data_io_write_ready;
  wire[127:0] data_io_resp_0;
  wire readArb_io_in_3_ready;
  wire readArb_io_in_2_ready;
  wire readArb_io_in_1_ready;
  wire readArb_io_out_valid;
  wire readArb_io_out_bits_way_en;
  wire[11:0] readArb_io_out_bits_addr;
  wire writeArb_io_in_1_ready;
  wire writeArb_io_out_valid;
  wire writeArb_io_out_bits_way_en;
  wire[11:0] writeArb_io_out_bits_addr;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[127:0] writeArb_io_out_bits_data;
  wire[63:0] amoalu_io_out;
  wire releaseArb_io_in_1_ready;
  wire releaseArb_io_in_0_ready;
  wire releaseArb_io_out_valid;
  wire[25:0] releaseArb_io_out_bits_addr;
  wire[1:0] releaseArb_io_out_bits_client_xact_id;
  wire[2:0] releaseArb_io_out_bits_master_xact_id;
  wire[511:0] releaseArb_io_out_bits_data;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire FlowThroughSerializer_0_io_in_ready;
  wire FlowThroughSerializer_0_io_out_valid;
  wire[1:0] FlowThroughSerializer_0_io_out_bits_header_src;
  wire[1:0] FlowThroughSerializer_0_io_out_bits_header_dst;
  wire[511:0] FlowThroughSerializer_0_io_out_bits_payload_data;
  wire[1:0] FlowThroughSerializer_0_io_out_bits_payload_client_xact_id;
  wire[2:0] FlowThroughSerializer_0_io_out_bits_payload_master_xact_id;
  wire[3:0] FlowThroughSerializer_0_io_out_bits_payload_g_type;
  wire wbArb_io_in_1_ready;
  wire wbArb_io_in_0_ready;
  wire wbArb_io_out_valid;
  wire[19:0] wbArb_io_out_bits_tag;
  wire[5:0] wbArb_io_out_bits_idx;
  wire wbArb_io_out_bits_way_en;
  wire[1:0] wbArb_io_out_bits_client_xact_id;
  wire[2:0] wbArb_io_out_bits_master_xact_id;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire dtlb_io_req_ready;
  wire dtlb_io_resp_miss;
  wire[18:0] dtlb_io_resp_ppn;
  wire dtlb_io_resp_xcpt_ld;
  wire dtlb_io_resp_xcpt_st;
  wire dtlb_io_ptw_req_valid;
  wire[29:0] dtlb_io_ptw_req_bits;
  wire mshrs_io_req_ready;
  wire mshrs_io_secondary_miss;
  wire mshrs_io_mem_req_valid;
  wire[25:0] mshrs_io_mem_req_bits_addr;
  wire[1:0] mshrs_io_mem_req_bits_client_xact_id;
  wire[511:0] mshrs_io_mem_req_bits_data;
  wire[2:0] mshrs_io_mem_req_bits_a_type;
  wire[5:0] mshrs_io_mem_req_bits_write_mask;
  wire[2:0] mshrs_io_mem_req_bits_subword_addr;
  wire[3:0] mshrs_io_mem_req_bits_atomic_opcode;
  wire mshrs_io_mem_resp_way_en;
  wire[11:0] mshrs_io_mem_resp_addr;
  wire mshrs_io_meta_read_valid;
  wire[5:0] mshrs_io_meta_read_bits_idx;
  wire mshrs_io_meta_write_valid;
  wire[5:0] mshrs_io_meta_write_bits_idx;
  wire mshrs_io_meta_write_bits_way_en;
  wire[19:0] mshrs_io_meta_write_bits_data_tag;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire mshrs_io_replay_valid;
  wire mshrs_io_replay_bits_kill;
  wire[2:0] mshrs_io_replay_bits_typ;
  wire mshrs_io_replay_bits_phys;
  wire[43:0] mshrs_io_replay_bits_addr;
  wire[63:0] mshrs_io_replay_bits_data;
  wire[7:0] mshrs_io_replay_bits_tag;
  wire[4:0] mshrs_io_replay_bits_cmd;
  wire mshrs_io_mem_finish_valid;
  wire[1:0] mshrs_io_mem_finish_bits_header_src;
  wire[1:0] mshrs_io_mem_finish_bits_header_dst;
  wire[2:0] mshrs_io_mem_finish_bits_payload_master_xact_id;
  wire mshrs_io_wb_req_valid;
  wire[19:0] mshrs_io_wb_req_bits_tag;
  wire[5:0] mshrs_io_wb_req_bits_idx;
  wire mshrs_io_wb_req_bits_way_en;
  wire[1:0] mshrs_io_wb_req_bits_client_xact_id;
  wire[2:0] mshrs_io_wb_req_bits_master_xact_id;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire mshrs_io_probe_rdy;
  wire mshrs_io_fence_rdy;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s2_recycle_next = {1{$random}};
    s1_valid = {1{$random}};
    s2_req_addr = {2{$random}};
    s1_req_addr = {2{$random}};
    s2_hit_state_state = {1{$random}};
    s2_tag_match_way = {1{$random}};
    R87 = {1{$random}};
    s2_valid = {1{$random}};
    s1_clk_en = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R191 = {2{$random}};
    R196 = {2{$random}};
    s2_store_bypass_data = {2{$random}};
    s4_req_data = {2{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_data = {2{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    R416 = {1{$random}};
    s2_repl_meta_coh_state = {1{$random}};
    s2_repl_meta_tag = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    block_miss = {1{$random}};
  end
`endif

  assign T367 = writeArb_io_in_1_ready | T368;
  assign T368 = T369 ^ 1'h1;
  assign T369 = T371 | T370;
  assign T370 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 4'h2;
  assign T371 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 4'h1;
  assign T372 = io_mem_release_ready;
  assign T161 = T168 ? s1_req_data : T162;
  assign T162 = T164 ? T163 : s2_req_data;
  assign T163 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T343 = reset ? 1'h0 : T26;
  assign T26 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T164 = s1_clk_en & s1_write;
  assign s1_write = T122 | T119;
  assign T119 = T121 | T120;
  assign T120 = s1_req_cmd == 5'h4;
  assign T19 = s2_recycle ? s2_req_cmd : T20;
  assign T20 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T21;
  assign T21 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T18 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T22;
  assign T22 = s2_recycle_ecc | s2_recycle_next;
  assign T342 = reset ? 1'h0 : T23;
  assign T23 = T28 ? T24 : s2_recycle_next;
  assign T24 = T25 & s2_recycle_ecc;
  assign T25 = s1_valid | s1_replay;
  assign T344 = reset ? 1'h0 : T27;
  assign T27 = io_cpu_req_ready & io_cpu_req_valid;
  assign T28 = s1_valid | s1_replay;
  assign s2_recycle_ecc = T46 & s2_data_correctable;
  assign s2_data_correctable = T44 & T29;
  assign T29 = T30 - 1'h1;
  assign T30 = 1'h1 << T31;
  assign T31 = T32 + 1'h1;
  assign T32 = s2_word_idx - s2_word_idx;
  assign s2_word_idx = s2_req_addr[2'h3:2'h3];
  assign T33 = s1_clk_en ? T345 : s2_req_addr;
  assign T345 = {12'h0, s1_addr};
  assign s1_addr = {dtlb_io_resp_ppn, T34};
  assign T34 = s1_req_addr[4'hc:1'h0];
  assign T35 = s2_recycle ? s2_req_addr : T36;
  assign T36 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T37;
  assign T37 = prober_io_meta_read_valid ? T347 : T38;
  assign T38 = wb_io_meta_read_valid ? T346 : T39;
  assign T39 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T346 = {12'h0, T40};
  assign T40 = T41 << 3'h6;
  assign T41 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T347 = {12'h0, T42};
  assign T42 = T43 << 3'h6;
  assign T43 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T44 = T45 >> s2_word_idx;
  assign T45 = 2'h0;
  assign T46 = T85 & s2_hit;
  assign s2_hit = T58 & T47;
  assign T47 = s2_hit_state_state == T48;
  assign T48 = T49;
  assign T49 = T50 ? 2'h3 : s2_hit_state_state;
  assign T50 = T54 | T51;
  assign T51 = T53 | T52;
  assign T52 = s2_req_cmd == 5'h4;
  assign T53 = s2_req_cmd[2'h3:2'h3];
  assign T54 = T56 | T55;
  assign T55 = s2_req_cmd == 5'h7;
  assign T56 = s2_req_cmd == 5'h1;
  assign T57 = s1_clk_en ? meta_io_resp_0_coh_state : s2_hit_state_state;
  assign T58 = s2_tag_match & T59;
  assign T59 = T68 ? T65 : T60;
  assign T60 = T62 | T61;
  assign T61 = s2_hit_state_state == 2'h3;
  assign T62 = T64 | T63;
  assign T63 = s2_hit_state_state == 2'h2;
  assign T64 = s2_hit_state_state == 2'h1;
  assign T65 = T67 | T66;
  assign T66 = s2_hit_state_state == 2'h3;
  assign T67 = s2_hit_state_state == 2'h2;
  assign T68 = T70 | T69;
  assign T69 = s2_req_cmd == 5'h6;
  assign T70 = T72 | T71;
  assign T71 = s2_req_cmd == 5'h3;
  assign T72 = T76 | T73;
  assign T73 = T75 | T74;
  assign T74 = s2_req_cmd == 5'h4;
  assign T75 = s2_req_cmd[2'h3:2'h3];
  assign T76 = T78 | T77;
  assign T77 = s2_req_cmd == 5'h7;
  assign T78 = s2_req_cmd == 5'h1;
  assign s2_tag_match = s2_tag_match_way != 1'h0;
  assign T79 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T80;
  assign T80 = T82 & T81;
  assign T81 = meta_io_resp_0_coh_state != 2'h0;
  assign T82 = s1_tag_eq_way;
  assign s1_tag_eq_way = T83;
  assign T83 = meta_io_resp_0_tag == T84;
  assign T84 = s1_addr >> 4'hc;
  assign T85 = s2_valid | s2_replay;
  assign s2_replay = R87 & T86;
  assign T86 = s2_req_cmd != 5'h5;
  assign T348 = reset ? 1'h0 : s1_replay;
  assign T349 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T88;
  assign T88 = io_cpu_req_bits_kill ^ 1'h1;
  assign T121 = s1_req_cmd[2'h3:2'h3];
  assign T122 = T124 | T123;
  assign T123 = s1_req_cmd == 5'h7;
  assign T124 = s1_req_cmd == 5'h1;
  assign T165 = s2_recycle ? s2_req_data : T166;
  assign T166 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T167;
  assign T167 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T168 = s1_clk_en & s1_recycled;
  assign T169 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T373 = s2_data_word[6'h3f:1'h0];
  assign s2_data_word = s2_store_bypass ? T354 : s2_data_word_prebypass;
  assign s2_data_word_prebypass = s2_data_uncorrected >> T186;
  assign T186 = {s2_word_idx, 6'h0};
  assign s2_data_uncorrected = T187;
  assign T187 = {T199, T188};
  assign T188 = s2_data_0[6'h3f:1'h0];
  assign s2_data_0 = T189;
  assign T189 = T190;
  assign T190 = {R196, R191};
  assign T352 = T192[6'h3f:1'h0];
  assign T192 = T194 ? T193 : T353;
  assign T353 = {64'h0, R191};
  assign T193 = data_io_resp_0 >> 1'h0;
  assign T194 = s1_clk_en & T195;
  assign T195 = s1_tag_eq_way;
  assign T197 = T194 ? T198 : R196;
  assign T198 = data_io_resp_0 >> 7'h40;
  assign T199 = s2_data_0[7'h7f:7'h40];
  assign T354 = {64'h0, s2_store_bypass_data};
  assign T200 = T260 ? T201 : s2_store_bypass_data;
  assign T201 = T245 ? amoalu_io_out : T202;
  assign T202 = T231 ? s3_req_data : s4_req_data;
  assign T203 = T204 ? s3_req_data : s4_req_data;
  assign T204 = s3_valid & metaReadArb_io_out_valid;
  assign T355 = reset ? 1'h0 : T205;
  assign T205 = T213 & T206;
  assign T206 = T210 | T207;
  assign T207 = T209 | T208;
  assign T208 = s2_req_cmd == 5'h4;
  assign T209 = s2_req_cmd[2'h3:2'h3];
  assign T210 = T212 | T211;
  assign T211 = s2_req_cmd == 5'h7;
  assign T212 = s2_req_cmd == 5'h1;
  assign T213 = T215 & T214;
  assign T214 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T171;
  assign T171 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = lrsc_valid & T172;
  assign T172 = lrsc_addr == T173;
  assign T173 = s2_req_addr >> 3'h6;
  assign T174 = T17 ? T175 : lrsc_addr;
  assign T175 = s2_req_addr >> 3'h6;
  assign T17 = T89 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T89 = T90 | s2_replay;
  assign T90 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T91;
  assign T91 = s2_valid & T92;
  assign T92 = s2_nack ^ 1'h1;
  assign s2_nack = T95 | s2_nack_miss;
  assign s2_nack_miss = T94 & T93;
  assign T93 = mshrs_io_req_ready ^ 1'h1;
  assign T94 = s2_hit ^ 1'h1;
  assign T95 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T96 = T102 ? s1_nack : s2_nack_hit;
  assign s1_nack = T101 | T97;
  assign T97 = T99 & T98;
  assign T98 = prober_io_req_ready ^ 1'h1;
  assign T99 = T100 == prober_io_meta_write_bits_idx;
  assign T100 = s1_req_addr[4'hb:3'h6];
  assign T101 = T405 & dtlb_io_resp_miss;
  assign T102 = s1_valid | s1_replay;
  assign lrsc_valid = lrsc_count != 5'h0;
  assign T341 = reset ? 5'h0 : T10;
  assign T10 = io_cpu_ptw_sret ? 5'h0 : T11;
  assign T11 = T103 ? 5'h0 : T12;
  assign T12 = T15 ? 5'h1f : T13;
  assign T13 = lrsc_valid ? T14 : lrsc_count;
  assign T14 = lrsc_count - 5'h1;
  assign T15 = T17 & T16;
  assign T16 = lrsc_valid ^ 1'h1;
  assign T103 = T89 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T215 = T216 | s2_replay;
  assign T216 = s2_valid_masked & s2_hit;
  assign T356 = T217[6'h3f:1'h0];
  assign T217 = T221 ? T219 : T357;
  assign T357 = {64'h0, T218};
  assign T218 = T221 ? s2_req_data : s3_req_data;
  assign T219 = s2_data_correctable ? s2_data_corrected : T358;
  assign T358 = {64'h0, amoalu_io_out};
  assign s2_data_corrected = T220;
  assign T220 = {T199, T188};
  assign T221 = T230 & T222;
  assign T222 = T223 | s2_data_correctable;
  assign T223 = T227 | T224;
  assign T224 = T226 | T225;
  assign T225 = s2_req_cmd == 5'h4;
  assign T226 = s2_req_cmd[2'h3:2'h3];
  assign T227 = T229 | T228;
  assign T228 = s2_req_cmd == 5'h7;
  assign T229 = s2_req_cmd == 5'h1;
  assign T230 = s2_valid | s2_replay;
  assign T231 = T240 & T232;
  assign T232 = T237 | T233;
  assign T233 = T236 | T234;
  assign T234 = s3_req_cmd == 5'h4;
  assign T235 = T221 ? s2_req_cmd : s3_req_cmd;
  assign T236 = s3_req_cmd[2'h3:2'h3];
  assign T237 = T239 | T238;
  assign T238 = s3_req_cmd == 5'h7;
  assign T239 = s3_req_cmd == 5'h1;
  assign T240 = s3_valid & T241;
  assign T241 = T359 == T242;
  assign T242 = s3_req_addr >> 2'h3;
  assign T243 = T221 ? s2_req_addr : s3_req_addr;
  assign T359 = {12'h0, T244};
  assign T244 = s1_addr >> 2'h3;
  assign T245 = T253 & T246;
  assign T246 = T250 | T247;
  assign T247 = T249 | T248;
  assign T248 = s2_req_cmd == 5'h4;
  assign T249 = s2_req_cmd[2'h3:2'h3];
  assign T250 = T252 | T251;
  assign T251 = s2_req_cmd == 5'h7;
  assign T252 = s2_req_cmd == 5'h1;
  assign T253 = T257 & T254;
  assign T254 = T360 == T255;
  assign T255 = s2_req_addr >> 2'h3;
  assign T360 = {12'h0, T256};
  assign T256 = s1_addr >> 2'h3;
  assign T257 = T259 & T258;
  assign T258 = s2_sc_fail ^ 1'h1;
  assign T259 = s2_valid_masked | s2_replay;
  assign T260 = s1_clk_en & T261;
  assign T261 = T276 | T262;
  assign T262 = T271 & T263;
  assign T263 = T268 | T264;
  assign T264 = T267 | T265;
  assign T265 = s4_req_cmd == 5'h4;
  assign T266 = T204 ? s3_req_cmd : s4_req_cmd;
  assign T267 = s4_req_cmd[2'h3:2'h3];
  assign T268 = T270 | T269;
  assign T269 = s4_req_cmd == 5'h7;
  assign T270 = s4_req_cmd == 5'h1;
  assign T271 = s4_valid & T272;
  assign T272 = T361 == T273;
  assign T273 = s4_req_addr >> 2'h3;
  assign T274 = T204 ? s3_req_addr : s4_req_addr;
  assign T361 = {12'h0, T275};
  assign T275 = s1_addr >> 2'h3;
  assign T362 = reset ? 1'h0 : s3_valid;
  assign T276 = T245 | T231;
  assign T277 = T260 ? 1'h1 : T278;
  assign T278 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T140 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T137 = s2_recycle ? s2_req_typ : T138;
  assign T138 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T139;
  assign T139 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T374 = s2_req_cmd[2'h3:1'h0];
  assign T375 = s2_req_addr[3'h5:1'h0];
  assign T376 = {s3_req_data, s3_req_data};
  assign T377 = 1'h1 << T378;
  assign T378 = T379;
  assign T379 = s3_req_addr[2'h3:2'h3];
  assign T380 = s3_req_addr[4'hb:1'h0];
  assign T381 = T221 ? s2_tag_match_way : s3_way;
  assign T382 = FlowThroughSerializer_0_io_out_bits_payload_data[7'h7f:1'h0];
  assign T383 = FlowThroughSerializer_0_io_out_valid & T384;
  assign T384 = T386 | T385;
  assign T385 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 4'h2;
  assign T386 = FlowThroughSerializer_0_io_out_bits_payload_g_type == 4'h1;
  assign T387 = T388 | T367;
  assign T388 = FlowThroughSerializer_0_io_out_valid ^ 1'h1;
  assign T389 = s2_req_addr[4'hb:1'h0];
  assign T390 = mshrs_io_replay_bits_addr[4'hb:1'h0];
  assign T391 = io_cpu_req_bits_addr[4'hb:1'h0];
  assign T392 = T393;
  assign T393 = {wdata_encoded_1, wdata_encoded_0};
  assign wdata_encoded_0 = writeArb_io_out_bits_data[6'h3f:1'h0];
  assign wdata_encoded_1 = writeArb_io_out_bits_data[7'h7f:7'h40];
  assign T394 = T395[3'h5:1'h0];
  assign T395 = s2_req_addr >> 3'h6;
  assign T396 = T397[3'h5:1'h0];
  assign T397 = io_cpu_req_bits_addr >> 3'h6;
  assign T398 = s2_recycle ? s2_req_phys : T399;
  assign T399 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T400;
  assign T400 = prober_io_meta_read_valid ? 1'h1 : T401;
  assign T401 = wb_io_meta_read_valid ? 1'h1 : T402;
  assign T402 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T403 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T404 = s1_req_addr >> 4'hd;
  assign T405 = T407 & T406;
  assign T406 = s1_req_phys ^ 1'h1;
  assign T407 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T411 | T408;
  assign T408 = T410 | T409;
  assign T409 = s1_req_cmd == 5'h3;
  assign T410 = s1_req_cmd == 5'h2;
  assign T411 = s1_read | s1_write;
  assign s1_read = T129 | T126;
  assign T126 = T128 | T127;
  assign T127 = s1_req_cmd == 5'h4;
  assign T128 = s1_req_cmd[2'h3:2'h3];
  assign T129 = T131 | T130;
  assign T130 = s1_req_cmd == 5'h6;
  assign T131 = s1_req_cmd == 5'h0;
  assign T412 = T367 & FlowThroughSerializer_0_io_out_valid;
  assign T413 = io_mem_acquire_ready;
  assign T414 = T415[1'h0:1'h0];
  assign T415 = s2_tag_match ? T418 : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R416;
  assign T417 = s1_clk_en ? 1'h0 : R416;
  assign T418 = {1'h0, s2_tag_match_way};
  assign T419 = s2_tag_match ? T421 : s2_repl_meta_coh_state;
  assign T420 = s1_clk_en ? meta_io_resp_0_coh_state : s2_repl_meta_coh_state;
  assign T421 = s2_hit_state_state;
  assign T422 = s2_tag_match ? T424 : s2_repl_meta_tag;
  assign T423 = s1_clk_en ? meta_io_resp_0_tag : s2_repl_meta_tag;
  assign T424 = s2_repl_meta_tag;
  assign T158 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T155 = s2_recycle ? s2_req_tag : T156;
  assign T156 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T157;
  assign T157 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T425 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T426 = s2_recycle ? s2_req_kill : T427;
  assign T427 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T428;
  assign T428 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T429 = s2_nack_hit ? 1'h0 : T430;
  assign T430 = T450 & T431;
  assign T431 = T439 | T432;
  assign T432 = T436 | T433;
  assign T433 = T435 | T434;
  assign T434 = s2_req_cmd == 5'h4;
  assign T435 = s2_req_cmd[2'h3:2'h3];
  assign T436 = T438 | T437;
  assign T437 = s2_req_cmd == 5'h7;
  assign T438 = s2_req_cmd == 5'h1;
  assign T439 = T447 | T440;
  assign T440 = T444 | T441;
  assign T441 = T443 | T442;
  assign T442 = s2_req_cmd == 5'h4;
  assign T443 = s2_req_cmd[2'h3:2'h3];
  assign T444 = T446 | T445;
  assign T445 = s2_req_cmd == 5'h6;
  assign T446 = s2_req_cmd == 5'h0;
  assign T447 = T449 | T448;
  assign T448 = s2_req_cmd == 5'h3;
  assign T449 = s2_req_cmd == 5'h2;
  assign T450 = s2_valid_masked & T451;
  assign T451 = s2_hit ^ 1'h1;
  assign probe_bits_p_type = io_mem_probe_bits_payload_p_type;
  assign probe_bits_master_xact_id = io_mem_probe_bits_payload_master_xact_id;
  assign probe_bits_addr = io_mem_probe_bits_payload_addr;
  assign T452 = probe_valid & T453;
  assign T453 = lrsc_valid ^ 1'h1;
  assign probe_valid = io_mem_probe_valid;
  assign io_mem_release_bits_payload_r_type = T0;
  assign T0 = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_payload_data = T1;
  assign T1 = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_payload_master_xact_id = T2;
  assign T2 = releaseArb_io_out_bits_master_xact_id;
  assign io_mem_release_bits_payload_client_xact_id = T3;
  assign T3 = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_payload_addr = T4;
  assign T4 = releaseArb_io_out_bits_addr;
  assign io_mem_release_bits_header_dst = T5;
  assign T5 = 2'h0;
  assign io_mem_release_bits_header_src = T6;
  assign T6 = 2'h0;
  assign io_mem_release_valid = T7;
  assign T7 = releaseArb_io_out_valid;
  assign io_mem_probe_ready = probe_ready;
  assign probe_ready = T8;
  assign T8 = prober_io_req_ready & T9;
  assign T9 = lrsc_valid ^ 1'h1;
  assign io_mem_finish_bits_payload_master_xact_id = mshrs_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mshrs_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = mshrs_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = mshrs_io_mem_finish_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_0_io_in_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = T104;
  assign T104 = mshrs_io_mem_req_bits_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = T105;
  assign T105 = mshrs_io_mem_req_bits_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = T106;
  assign T106 = mshrs_io_mem_req_bits_write_mask;
  assign io_mem_acquire_bits_payload_a_type = T107;
  assign T107 = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_payload_data = T108;
  assign T108 = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_payload_client_xact_id = T109;
  assign T109 = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = T110;
  assign T110 = mshrs_io_mem_req_bits_addr;
  assign io_mem_acquire_bits_header_dst = T111;
  assign T111 = 2'h0;
  assign io_mem_acquire_bits_header_src = T112;
  assign T112 = 2'h0;
  assign io_mem_acquire_valid = T113;
  assign T113 = mshrs_io_mem_req_valid;
  assign io_cpu_ordered = T114;
  assign T114 = T116 & T115;
  assign T115 = s2_valid ^ 1'h1;
  assign T116 = mshrs_io_fence_rdy & T117;
  assign T117 = s1_valid ^ 1'h1;
  assign io_cpu_ptw_req_bits = dtlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_xcpt_pf_st = T118;
  assign T118 = s1_write & dtlb_io_resp_xcpt_st;
  assign io_cpu_xcpt_pf_ld = T125;
  assign T125 = s1_read & dtlb_io_resp_xcpt_ld;
  assign io_cpu_xcpt_ma_st = T132;
  assign T132 = s1_write & misaligned;
  assign misaligned = T141 | T133;
  assign T133 = T136 & T134;
  assign T134 = T135 != 3'h0;
  assign T135 = s1_req_addr[2'h2:1'h0];
  assign T136 = s1_req_typ == 3'h3;
  assign T141 = T148 | T142;
  assign T142 = T145 & T143;
  assign T143 = T144 != 2'h0;
  assign T144 = s1_req_addr[1'h1:1'h0];
  assign T145 = T147 | T146;
  assign T146 = s1_req_typ == 3'h6;
  assign T147 = s1_req_typ == 3'h2;
  assign T148 = T151 & T149;
  assign T149 = T150 != 1'h0;
  assign T150 = s1_req_addr[1'h0:1'h0];
  assign T151 = T153 | T152;
  assign T152 = s1_req_typ == 3'h5;
  assign T153 = s1_req_typ == 3'h1;
  assign io_cpu_xcpt_ma_ld = T154;
  assign T154 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T159;
  assign T159 = s1_replay & T160;
  assign T160 = s1_read | s1_sc;
  assign s1_sc = s1_req_cmd == 5'h7;
  assign io_cpu_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_bits_cmd = T350;
  assign T350 = s2_req_cmd[2'h3:1'h0];
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_data_subword = T170;
  assign T170 = T176 | T351;
  assign T351 = {63'h0, s2_sc_fail};
  assign T176 = {T308, T177};
  assign T177 = s2_sc ? 8'h0 : T178;
  assign T178 = T307 ? T306 : T179;
  assign T179 = T180[3'h7:1'h0];
  assign T180 = {T298, T181};
  assign T181 = T297 ? T296 : T182;
  assign T182 = T183[4'hf:1'h0];
  assign T183 = {T281, T184};
  assign T184 = T280 ? T279 : T185;
  assign T185 = s2_data_word[5'h1f:1'h0];
  assign T279 = s2_data_word[6'h3f:6'h20];
  assign T280 = s2_req_addr[2'h2:2'h2];
  assign T281 = T293 ? T283 : T282;
  assign T282 = s2_data_word[6'h3f:6'h20];
  assign T283 = 32'h0 - T363;
  assign T363 = {31'h0, T284};
  assign T284 = T286 & T285;
  assign T285 = T184[5'h1f:5'h1f];
  assign T286 = T288 | T287;
  assign T287 = s2_req_typ == 3'h3;
  assign T288 = T290 | T289;
  assign T289 = s2_req_typ == 3'h2;
  assign T290 = T292 | T291;
  assign T291 = s2_req_typ == 3'h1;
  assign T292 = s2_req_typ == 3'h0;
  assign T293 = T295 | T294;
  assign T294 = s2_req_typ == 3'h6;
  assign T295 = s2_req_typ == 3'h2;
  assign T296 = T183[5'h1f:5'h10];
  assign T297 = s2_req_addr[1'h1:1'h1];
  assign T298 = T303 ? T300 : T299;
  assign T299 = T183[6'h3f:5'h10];
  assign T300 = 48'h0 - T364;
  assign T364 = {47'h0, T301};
  assign T301 = T286 & T302;
  assign T302 = T181[4'hf:4'hf];
  assign T303 = T305 | T304;
  assign T304 = s2_req_typ == 3'h5;
  assign T305 = s2_req_typ == 3'h1;
  assign T306 = T180[4'hf:4'h8];
  assign T307 = s2_req_addr[1'h0:1'h0];
  assign T308 = T313 ? T310 : T309;
  assign T309 = T180[6'h3f:4'h8];
  assign T310 = 56'h0 - T365;
  assign T365 = {55'h0, T311};
  assign T311 = T286 & T312;
  assign T312 = T177[3'h7:3'h7];
  assign T313 = s2_sc | T314;
  assign T314 = T316 | T315;
  assign T315 = s2_req_typ == 3'h4;
  assign T316 = s2_req_typ == 3'h0;
  assign io_cpu_resp_bits_data = T183;
  assign io_cpu_resp_bits_has_data = T317;
  assign T317 = T318 | s2_sc;
  assign T318 = T322 | T319;
  assign T319 = T321 | T320;
  assign T320 = s2_req_cmd == 5'h4;
  assign T321 = s2_req_cmd[2'h3:2'h3];
  assign T322 = T324 | T323;
  assign T323 = s2_req_cmd == 5'h6;
  assign T324 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T325;
  assign T325 = s2_valid & s2_nack;
  assign io_cpu_resp_valid = T326;
  assign T326 = T328 & T327;
  assign T327 = s2_data_correctable ^ 1'h1;
  assign T328 = s2_replay | T329;
  assign T329 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T330;
  assign T330 = block_miss ? 1'h0 : T331;
  assign T331 = T338 ? 1'h0 : T332;
  assign T332 = T337 ? 1'h0 : T333;
  assign T333 = T334 == 1'h0;
  assign T334 = T336 & T335;
  assign T335 = io_cpu_req_bits_phys ^ 1'h1;
  assign T336 = dtlb_io_req_ready ^ 1'h1;
  assign T337 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T338 = readArb_io_in_3_ready ^ 1'h1;
  assign T366 = reset ? 1'h0 : T339;
  assign T339 = T340 & s2_nack_miss;
  assign T340 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_tag( wbArb_io_out_bits_tag ),
       .io_req_bits_idx( wbArb_io_out_bits_idx ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_master_xact_id( wbArb_io_out_bits_master_xact_id ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( s2_data_corrected ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr( wb_io_release_bits_addr ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_master_xact_id( wb_io_release_bits_master_xact_id ),
       .io_release_bits_data( wb_io_release_bits_data ),
       .io_release_bits_r_type( wb_io_release_bits_r_type )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T452 ),
       .io_req_bits_addr( probe_bits_addr ),
       .io_req_bits_master_xact_id( probe_bits_master_xact_id ),
       .io_req_bits_p_type( probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr( prober_io_rep_bits_addr ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_master_xact_id( prober_io_rep_bits_master_xact_id ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_tag( prober_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( prober_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( prober_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_line_state_state( s2_hit_state_state )
  );
  `ifndef SYNTHESIS
    assign prober.io_req_bits_client_xact_id = {1{$random}};
  `endif
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T429 ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_data( s2_req_data ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_tag_match( s2_tag_match ),
       .io_req_bits_old_meta_tag( T422 ),
       .io_req_bits_old_meta_coh_state( T419 ),
       .io_req_bits_way_en( T414 ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( T413 ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr( mshrs_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_write_mask( mshrs_io_mem_req_bits_write_mask ),
       .io_mem_req_bits_subword_addr( mshrs_io_mem_req_bits_subword_addr ),
       .io_mem_req_bits_atomic_opcode( mshrs_io_mem_req_bits_atomic_opcode ),
       .io_mem_resp_way_en( mshrs_io_mem_resp_way_en ),
       .io_mem_resp_addr( mshrs_io_mem_resp_addr ),
       //.io_mem_resp_wmask(  )
       //.io_mem_resp_data(  )
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       //.io_replay_bits_sdq_id(  )
       .io_mem_grant_valid( T412 ),
       .io_mem_grant_bits_header_src( FlowThroughSerializer_0_io_out_bits_header_src ),
       .io_mem_grant_bits_header_dst( FlowThroughSerializer_0_io_out_bits_header_dst ),
       .io_mem_grant_bits_payload_data( FlowThroughSerializer_0_io_out_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( FlowThroughSerializer_0_io_out_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( FlowThroughSerializer_0_io_out_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( FlowThroughSerializer_0_io_out_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( mshrs_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( mshrs_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( mshrs_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( mshrs_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( mshrs_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T405 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T404 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_resp_miss( dtlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits( dtlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state )
  );
  Arbiter_0 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T396 ),
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T394 ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx )
       //.io_chosen(  )
  );
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T392 ),
       .io_resp_0( data_io_resp_0 )
  );
  Arbiter_2 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 1'h1 ),
       .io_in_3_bits_addr( T391 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 1'h1 ),
       .io_in_1_bits_addr( T390 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 1'h1 ),
       .io_in_0_bits_addr( T389 ),
       .io_out_ready( T387 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_3 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T383 ),
       .io_in_1_bits_way_en( mshrs_io_mem_resp_way_en ),
       .io_in_1_bits_addr( mshrs_io_mem_resp_addr ),
       .io_in_1_bits_wmask( 2'h3 ),
       .io_in_1_bits_data( T382 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T380 ),
       .io_in_0_bits_wmask( T377 ),
       .io_in_0_bits_data( T376 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T375 ),
       .io_cmd( T374 ),
       .io_typ( s2_req_typ ),
       .io_lhs( T373 ),
       .io_rhs( s2_req_data ),
       .io_out( amoalu_io_out )
  );
  Arbiter_4 releaseArb(
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr( prober_io_rep_bits_addr ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( prober_io_rep_bits_master_xact_id ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr( wb_io_release_bits_addr ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( wb_io_release_bits_master_xact_id ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_out_ready( T372 ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr( releaseArb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( releaseArb_io_out_bits_master_xact_id ),
       .io_out_bits_data( releaseArb_io_out_bits_data ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  FlowThroughSerializer_0 FlowThroughSerializer_0(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_0_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( T367 ),
       .io_out_valid( FlowThroughSerializer_0_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( FlowThroughSerializer_0_io_out_bits_header_dst ),
       .io_out_bits_payload_data( FlowThroughSerializer_0_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( FlowThroughSerializer_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_0_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_0_io_out_bits_payload_g_type )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_5 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( mshrs_io_wb_req_bits_master_xact_id ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_tag( prober_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( prober_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( prober_io_wb_req_bits_master_xact_id ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_tag( wbArb_io_out_bits_tag ),
       .io_out_bits_idx( wbArb_io_out_bits_idx ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( wbArb_io_out_bits_master_xact_id ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
    if(T168) begin
      s2_req_data <= s1_req_data;
    end else if(T164) begin
      s2_req_data <= T163;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T26;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T28) begin
      s2_recycle_next <= T24;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T27;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T345;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T347;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T346;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_hit_state_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(reset) begin
      R87 <= 1'h0;
    end else begin
      R87 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R191 <= T352;
    if(T194) begin
      R196 <= T198;
    end
    if(T260) begin
      s2_store_bypass_data <= T201;
    end
    if(T204) begin
      s4_req_data <= s3_req_data;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T205;
    end
    if(T17) begin
      lrsc_addr <= T175;
    end
    if(T102) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_ptw_sret) begin
      lrsc_count <= 5'h0;
    end else if(T103) begin
      lrsc_count <= 5'h0;
    end else if(T15) begin
      lrsc_count <= 5'h1f;
    end else if(lrsc_valid) begin
      lrsc_count <= T14;
    end
    s3_req_data <= T356;
    if(T221) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T221) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T204) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T204) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T260) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T221) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    if(s1_clk_en) begin
      R416 <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_repl_meta_coh_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_repl_meta_tag <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T339;
    end
  end
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [29:0] io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [29:0] io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output[29:0] io_out_bits,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T28;
  wire T6;
  wire T7;
  wire[29:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T28 = reset ? 1'h0 : T6;
  assign T6 = T7 ? T0 : R5;
  assign T7 = io_out_ready & io_out_valid;
  assign io_out_bits = T8;
  assign T8 = T9 ? io_in_1_bits : io_in_0_bits;
  assign T9 = T0;
  assign io_out_valid = T10;
  assign T10 = T9 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = T19 | T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = T17 | T15;
  assign T15 = io_in_1_valid & T16;
  assign T16 = R5 < 1'h1;
  assign T17 = io_in_0_valid & T18;
  assign T18 = R5 < 1'h0;
  assign T19 = R5 < 1'h0;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = T25 | T22;
  assign T22 = T23 ^ 1'h1;
  assign T23 = T24 | io_in_0_valid;
  assign T24 = T17 | T15;
  assign T25 = T27 & T26;
  assign T26 = R5 < 1'h1;
  assign T27 = T17 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T7) begin
      R5 <= T0;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [29:0] io_requestor_1_req_bits,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[18:0] io_requestor_1_resp_bits_ppn,
    output[5:0] io_requestor_1_resp_bits_perm,
    output[7:0] io_requestor_1_status_ip,
    output[7:0] io_requestor_1_status_im,
    output[6:0] io_requestor_1_status_zero,
    output io_requestor_1_status_er,
    output io_requestor_1_status_vm,
    output io_requestor_1_status_s64,
    output io_requestor_1_status_u64,
    output io_requestor_1_status_ef,
    output io_requestor_1_status_pei,
    output io_requestor_1_status_ei,
    output io_requestor_1_status_ps,
    output io_requestor_1_status_s,
    output io_requestor_1_invalidate,
    output io_requestor_1_sret,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [29:0] io_requestor_0_req_bits,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[18:0] io_requestor_0_resp_bits_ppn,
    output[5:0] io_requestor_0_resp_bits_perm,
    output[7:0] io_requestor_0_status_ip,
    output[7:0] io_requestor_0_status_im,
    output[6:0] io_requestor_0_status_zero,
    output io_requestor_0_status_er,
    output io_requestor_0_status_vm,
    output io_requestor_0_status_s64,
    output io_requestor_0_status_u64,
    output io_requestor_0_status_ef,
    output io_requestor_0_status_pei,
    output io_requestor_0_status_ei,
    output io_requestor_0_status_ps,
    output io_requestor_0_status_s,
    output io_requestor_0_invalidate,
    output io_requestor_0_sret,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    //output[63:0] io_mem_req_bits_data
    //output[7:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    input  io_mem_resp_valid,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    //input  io_mem_ptw_req_valid
    //input [29:0] io_mem_ptw_req_bits
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_sret,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s
);

  wire T79;
  reg [2:0] state;
  wire[2:0] T75;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T14;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T37;
  wire T38;
  wire T39;
  reg [1:0] count;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T36;
  wire T40;
  wire T34;
  wire T35;
  wire[43:0] T74;
  wire[31:0] T0;
  wire[28:0] T1;
  wire[28:0] T2;
  wire[9:0] vpn_idx;
  wire[9:0] T3;
  wire[9:0] T4;
  wire[9:0] T5;
  reg [29:0] r_req_vpn;
  wire[29:0] T6;
  wire T7;
  wire[9:0] T8;
  wire[19:0] T9;
  wire T10;
  wire[1:0] T11;
  wire[9:0] T41;
  wire[29:0] T42;
  wire T43;
  wire[18:0] T44;
  reg [63:0] r_pte;
  wire[63:0] T45;
  wire[63:0] T46;
  wire[63:0] T76;
  wire[31:0] T47;
  wire[12:0] T48;
  wire[18:0] T49;
  wire T50;
  wire[5:0] T51;
  wire[18:0] T77;
  wire[30:0] T52;
  wire[30:0] resp_ppn;
  wire[30:0] T53;
  wire[30:0] T54;
  wire[19:0] T55;
  wire[10:0] T56;
  wire[30:0] T57;
  wire[9:0] T58;
  wire[20:0] T59;
  wire T60;
  wire[1:0] T61;
  wire[30:0] r_resp_ppn;
  wire T62;
  wire resp_err;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  reg  r_req_dest;
  wire T67;
  wire resp_val;
  wire T68;
  wire T69;
  wire[5:0] T70;
  wire[18:0] T78;
  wire[30:0] T71;
  wire T72;
  wire T73;
  wire arb_io_in_1_ready;
  wire arb_io_in_0_ready;
  wire arb_io_out_valid;
  wire[29:0] arb_io_out_bits;
  wire arb_io_chosen;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    r_req_vpn = {1{$random}};
    r_pte = {2{$random}};
    r_req_dest = {1{$random}};
  end
`endif

  assign T79 = state == 3'h0;
  assign T75 = reset ? 3'h0 : T15;
  assign T15 = T35 ? 3'h0 : T16;
  assign T16 = T34 ? 3'h0 : T17;
  assign T17 = T37 ? 3'h1 : T18;
  assign T18 = T29 ? 3'h3 : T19;
  assign T19 = T28 ? 3'h4 : T20;
  assign T20 = T26 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h1 : state;
  assign T23 = T14 & arb_io_out_valid;
  assign T14 = 3'h0 == state;
  assign T24 = T25 & io_mem_req_ready;
  assign T25 = 3'h1 == state;
  assign T26 = T27 & io_mem_resp_bits_nack;
  assign T27 = 3'h2 == state;
  assign T28 = T27 & io_mem_resp_valid;
  assign T29 = T32 & T30;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_mem_resp_bits_data[1'h1:1'h1];
  assign T32 = T28 & T33;
  assign T33 = io_mem_resp_bits_data[1'h0:1'h0];
  assign T37 = T32 & T38;
  assign T38 = T40 & T39;
  assign T39 = count < 2'h2;
  assign T12 = T37 ? T36 : T13;
  assign T13 = T14 ? 2'h0 : count;
  assign T36 = count + 2'h1;
  assign T40 = T30 ^ 1'h1;
  assign T34 = 3'h3 == state;
  assign T35 = 3'h4 == state;
  assign io_mem_req_bits_cmd = 5'h0;
  assign io_mem_req_bits_addr = T74;
  assign T74 = {12'h0, T0};
  assign T0 = T1 << 2'h3;
  assign T1 = T2;
  assign T2 = {T44, vpn_idx};
  assign vpn_idx = T43 ? T41 : T3;
  assign T3 = T10 ? T8 : T4;
  assign T4 = T5[4'h9:1'h0];
  assign T5 = r_req_vpn >> 5'h14;
  assign T6 = T7 ? arb_io_out_bits : r_req_vpn;
  assign T7 = T79 & arb_io_out_valid;
  assign T8 = T9[4'h9:1'h0];
  assign T9 = r_req_vpn >> 4'ha;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = count;
  assign T41 = T42[4'h9:1'h0];
  assign T42 = r_req_vpn >> 1'h0;
  assign T43 = T11[1'h1:1'h1];
  assign T44 = r_pte[5'h1f:4'hd];
  assign T45 = io_mem_resp_valid ? io_mem_resp_bits_data : T46;
  assign T46 = T7 ? T76 : r_pte;
  assign T76 = {32'h0, T47};
  assign T47 = {T49, T48};
  assign T48 = io_mem_resp_bits_data[4'hc:1'h0];
  assign T49 = io_dpath_ptbr[5'h1f:4'hd];
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_valid = T50;
  assign T50 = state == 3'h1;
  assign io_requestor_0_sret = io_dpath_sret;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_s = io_dpath_status_s;
  assign io_requestor_0_status_ps = io_dpath_status_ps;
  assign io_requestor_0_status_ei = io_dpath_status_ei;
  assign io_requestor_0_status_pei = io_dpath_status_pei;
  assign io_requestor_0_status_ef = io_dpath_status_ef;
  assign io_requestor_0_status_u64 = io_dpath_status_u64;
  assign io_requestor_0_status_s64 = io_dpath_status_s64;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_er = io_dpath_status_er;
  assign io_requestor_0_status_zero = io_dpath_status_zero;
  assign io_requestor_0_status_im = io_dpath_status_im;
  assign io_requestor_0_status_ip = io_dpath_status_ip;
  assign io_requestor_0_resp_bits_perm = T51;
  assign T51 = r_pte[4'h8:2'h3];
  assign io_requestor_0_resp_bits_ppn = T77;
  assign T77 = T52[5'h12:1'h0];
  assign T52 = resp_ppn;
  assign resp_ppn = T62 ? r_resp_ppn : T53;
  assign T53 = T60 ? T57 : T54;
  assign T54 = {T56, T55};
  assign T55 = r_req_vpn[5'h13:1'h0];
  assign T56 = r_resp_ppn >> 5'h14;
  assign T57 = {T59, T58};
  assign T58 = r_req_vpn[4'h9:1'h0];
  assign T59 = r_resp_ppn >> 4'ha;
  assign T60 = T61[1'h0:1'h0];
  assign T61 = count;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hd;
  assign T62 = T61[1'h1:1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = T64 | T63;
  assign T63 = state == 3'h2;
  assign T64 = state == 3'h4;
  assign io_requestor_0_resp_valid = T65;
  assign T65 = resp_val & T66;
  assign T66 = r_req_dest == 1'h0;
  assign T67 = T7 ? arb_io_chosen : r_req_dest;
  assign resp_val = T69 | T68;
  assign T68 = state == 3'h4;
  assign T69 = state == 3'h3;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_sret = io_dpath_sret;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_s = io_dpath_status_s;
  assign io_requestor_1_status_ps = io_dpath_status_ps;
  assign io_requestor_1_status_ei = io_dpath_status_ei;
  assign io_requestor_1_status_pei = io_dpath_status_pei;
  assign io_requestor_1_status_ef = io_dpath_status_ef;
  assign io_requestor_1_status_u64 = io_dpath_status_u64;
  assign io_requestor_1_status_s64 = io_dpath_status_s64;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_er = io_dpath_status_er;
  assign io_requestor_1_status_zero = io_dpath_status_zero;
  assign io_requestor_1_status_im = io_dpath_status_im;
  assign io_requestor_1_status_ip = io_dpath_status_ip;
  assign io_requestor_1_resp_bits_perm = T70;
  assign T70 = r_pte[4'h8:2'h3];
  assign io_requestor_1_resp_bits_ppn = T78;
  assign T78 = T71[5'h12:1'h0];
  assign T71 = resp_ppn;
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T72;
  assign T72 = resp_val & T73;
  assign T73 = r_req_dest == 1'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  RRArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits( io_requestor_1_req_bits ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits( io_requestor_0_req_bits ),
       .io_out_ready( T79 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits( arb_io_out_bits ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h0;
    end else if(T37) begin
      state <= 3'h1;
    end else if(T29) begin
      state <= 3'h3;
    end else if(T28) begin
      state <= 3'h4;
    end else if(T26) begin
      state <= 3'h1;
    end else if(T24) begin
      state <= 3'h2;
    end else if(T23) begin
      state <= 3'h1;
    end
    if(T37) begin
      count <= T36;
    end else if(T14) begin
      count <= 2'h0;
    end
    if(T7) begin
      r_req_vpn <= arb_io_out_bits;
    end
    if(io_mem_resp_valid) begin
      r_pte <= io_mem_resp_bits_data;
    end else if(T7) begin
      r_pte <= T76;
    end
    if(T7) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module Control(input clk, input reset,
    output[2:0] io_dpath_sel_pc,
    output io_dpath_killd,
    output io_dpath_ren_1,
    output io_dpath_ren_0,
    output[2:0] io_dpath_sel_alu2,
    output[1:0] io_dpath_sel_alu1,
    output[2:0] io_dpath_sel_imm,
    output io_dpath_fn_dw,
    output[3:0] io_dpath_fn_alu,
    output io_dpath_div_mul_val,
    output io_dpath_div_mul_kill,
    //output io_dpath_div_val
    //output io_dpath_div_kill
    output[2:0] io_dpath_csr,
    output io_dpath_sret,
    output io_dpath_mem_load,
    output io_dpath_wb_load,
    output io_dpath_ex_fp_val,
    output io_dpath_mem_fp_val,
    output io_dpath_ex_wen,
    output io_dpath_ex_valid,
    output io_dpath_mem_jalr,
    output io_dpath_mem_branch,
    output io_dpath_mem_wen,
    output io_dpath_wb_wen,
    output[2:0] io_dpath_ex_mem_type,
    output io_dpath_ex_rs2_val,
    output io_dpath_ex_rocc_val,
    output io_dpath_mem_rocc_val,
    output io_dpath_bypass_1,
    output io_dpath_bypass_0,
    output[1:0] io_dpath_bypass_src_1,
    output[1:0] io_dpath_bypass_src_0,
    output io_dpath_ll_ready,
    output io_dpath_retire,
    output io_dpath_exception,
    output[63:0] io_dpath_cause,
    output io_dpath_badvaddr_wen,
    input [31:0] io_dpath_inst,
    //input  io_dpath_jalr_eq
    input  io_dpath_mem_br_taken,
    input  io_dpath_mem_misprediction,
    input  io_dpath_div_mul_rdy,
    input  io_dpath_ll_wen,
    input [4:0] io_dpath_ll_waddr,
    input [4:0] io_dpath_ex_waddr,
    input  io_dpath_mem_rs1_ra,
    input [4:0] io_dpath_mem_waddr,
    input [4:0] io_dpath_wb_waddr,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s,
    input  io_dpath_fp_sboard_clr,
    input [4:0] io_dpath_fp_sboard_clra,
    input  io_dpath_csr_replay,
    output io_imem_req_valid,
    //output[43:0] io_imem_req_bits_pc
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_index,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[2:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[3:0] io_imem_btb_update_bits_prediction_bits_bht_index,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    //output[42:0] io_imem_btb_update_bits_pc
    //output[42:0] io_imem_btb_update_bits_target
    //output[42:0] io_imem_btb_update_bits_returnAddr
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_incorrectTarget,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    //output[43:0] io_dmem_req_bits_addr
    //output[63:0] io_dmem_req_bits_data
    //output[7:0] io_dmem_req_bits_tag
    output[4:0] io_dmem_req_bits_cmd,
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output io_fpu_valid,
    //input  io_fpu_fcsr_rdy
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    //input [4:0] io_fpu_dec_cmd
    //input  io_fpu_dec_ldst
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    //input  io_fpu_dec_swap23
    //input  io_fpu_dec_single
    //input  io_fpu_dec_fromint
    //input  io_fpu_dec_toint
    //input  io_fpu_dec_fastpipe
    //input  io_fpu_dec_fma
    //input  io_fpu_dec_round
    //input  io_fpu_sboard_set
    //input  io_fpu_sboard_clr
    //input [4:0] io_fpu_sboard_clra
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire T0;
  reg  wb_reg_xcpt;
  wire T1;
  wire T2;
  wire take_pc_wb;
  wire T3;
  reg  wb_reg_sret;
  wire T4;
  wire T5;
  wire T6;
  reg  mem_reg_replay;
  wire T7;
  wire replay_ex;
  wire replay_ex_other;
  reg  mem_reg_replay_next;
  wire T8;
  reg  ex_reg_replay_next;
  wire T9;
  wire T10;
  wire id_csr_flush;
  wire T11;
  wire T12;
  wire T13;
  wire[11:0] T14;
  wire[11:0] id_csr_addr;
  wire T15;
  wire[11:0] T16;
  wire T17;
  wire id_csr_wen;
  wire T18;
  wire T19;
  wire T20;
  wire[1:0] id_csr;
  wire T21;
  wire[31:0] T22;
  wire T23;
  wire[31:0] T24;
  wire T25;
  wire T26;
  wire[4:0] id_raddr1;
  wire id_csr_en;
  wire id_replay_next;
  wire[31:0] T27;
  wire ctrl_killd;
  wire T28;
  wire ctrl_draind;
  wire id_interrupt;
  wire id_interrupt_unmasked;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire ctrl_stalld;
  wire id_do_fence;
  wire T60;
  wire T61;
  wire T62;
  wire id_mem_val;
  wire T63;
  wire[31:0] T64;
  wire T65;
  wire T66;
  wire[31:0] T67;
  wire T68;
  wire T69;
  wire[31:0] T70;
  wire T71;
  wire T72;
  wire[31:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T76;
  wire T77;
  wire[31:0] T78;
  reg  id_reg_fence;
  wire T665;
  wire T79;
  wire T80;
  wire id_fence_next;
  wire T81;
  wire id_amo_rl;
  wire id_amo;
  wire[31:0] T82;
  wire id_fence;
  wire[31:0] T83;
  wire T84;
  wire id_fence_i;
  wire[31:0] T85;
  wire T86;
  wire id_amo_aq;
  wire id_mem_busy;
  reg  ex_reg_mem_val;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire id_sboard_hazard;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[4:0] T98;
  wire[4:0] T99;
  wire[4:0] id_waddr;
  wire T100;
  wire[31:0] T101;
  wire[31:0] T102;
  wire[31:0] T103;
  wire[31:0] T104;
  reg [31:0] R105;
  wire[31:0] T666;
  wire[31:0] T106;
  wire[31:0] T107;
  wire[31:0] T108;
  wire[31:0] T109;
  wire[31:0] T110;
  wire T111;
  wire wb_set_sboard;
  reg  wb_reg_rocc_val;
  wire T112;
  reg  mem_reg_rocc_val;
  wire T113;
  reg  ex_reg_rocc_val;
  wire T114;
  wire T115;
  wire T116;
  wire wb_dcache_miss;
  wire T117;
  reg  wb_reg_mem_val;
  wire T118;
  reg  mem_reg_mem_val;
  wire T119;
  reg  wb_reg_div_mul_val;
  wire T120;
  reg  mem_reg_div_mul_val;
  wire T121;
  reg  ex_reg_div_mul_val;
  wire T122;
  wire T123;
  wire id_div_val;
  wire[31:0] T124;
  wire id_mul_val;
  wire[31:0] T125;
  wire T126;
  wire id_wen_not0;
  wire T127;
  wire id_wen;
  wire T128;
  wire[31:0] T129;
  wire T130;
  wire T131;
  wire[31:0] T132;
  wire T133;
  wire T134;
  wire[31:0] T135;
  wire T136;
  wire T137;
  wire[31:0] T138;
  wire T139;
  wire id_jal;
  wire[31:0] T140;
  wire T141;
  wire T142;
  wire[31:0] T143;
  wire T144;
  wire[31:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire[4:0] T152;
  wire[4:0] id_raddr2;
  wire T153;
  wire id_renx2_not0;
  wire T154;
  wire id_renx2;
  wire T155;
  wire[31:0] T156;
  wire T157;
  wire T158;
  wire[31:0] T159;
  wire T160;
  wire[31:0] T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire[4:0] T166;
  wire[4:0] T167;
  wire T168;
  wire id_renx1_not0;
  wire T169;
  wire id_renx1;
  wire T170;
  wire[31:0] T171;
  wire T172;
  wire T173;
  wire[31:0] T174;
  wire T175;
  wire T176;
  wire[31:0] T177;
  wire T178;
  wire T179;
  wire[31:0] T180;
  wire T181;
  wire[31:0] T182;
  wire T183;
  wire id_wb_hazard;
  wire T184;
  wire T185;
  reg  wb_reg_fp_val;
  wire T186;
  reg  mem_reg_fp_val;
  wire T187;
  reg  ex_reg_fp_val;
  wire T188;
  wire fp_data_hazard_wb;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire[4:0] id_raddr3;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  reg  wb_reg_fp_wen;
  wire T200;
  reg  mem_reg_fp_wen;
  wire T201;
  reg  ex_reg_fp_wen;
  wire T202;
  wire T203;
  wire data_hazard_wb;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  reg  wb_reg_wen;
  wire T212;
  reg  mem_reg_wen;
  wire T213;
  reg  ex_reg_wen;
  wire T214;
  wire T215;
  wire id_mem_hazard;
  wire T216;
  wire fp_data_hazard_mem;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  reg  mem_mem_cmd_bh;
  wire T234;
  wire ex_slow_bypass;
  wire T235;
  wire T236;
  reg [2:0] ex_reg_mem_type;
  wire[2:0] T237;
  wire[2:0] T238;
  wire[2:0] id_mem_type;
  wire[1:0] T239;
  wire T240;
  wire[31:0] T241;
  wire T242;
  wire[31:0] T243;
  wire T244;
  wire[31:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg [4:0] ex_reg_mem_cmd;
  wire[4:0] T253;
  wire[4:0] id_mem_cmd;
  wire[3:0] T254;
  wire[2:0] T255;
  wire[1:0] T256;
  wire T257;
  wire T258;
  wire[31:0] T259;
  wire T260;
  wire T261;
  wire[31:0] T262;
  wire T263;
  wire[31:0] T264;
  wire T265;
  wire T266;
  wire[31:0] T267;
  wire T268;
  wire[31:0] T269;
  wire T270;
  wire T271;
  wire[31:0] T272;
  wire T273;
  wire T274;
  wire[31:0] T275;
  wire T276;
  wire[31:0] T277;
  wire T278;
  wire T279;
  reg [1:0] mem_reg_csr;
  wire[1:0] T280;
  reg [1:0] ex_reg_csr;
  wire[1:0] T281;
  wire data_hazard_mem;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire id_ex_hazard;
  wire T290;
  wire T291;
  wire fp_data_hazard_ex;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  reg  ex_reg_jalr;
  wire T309;
  wire id_jalr;
  wire[31:0] T310;
  wire T311;
  wire data_hazard_ex;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire take_pc;
  wire take_pc_mem;
  wire T321;
  reg  mem_reg_jal;
  wire T322;
  reg  ex_reg_jal;
  wire T323;
  wire T324;
  reg  mem_reg_jalr;
  wire T325;
  reg  mem_reg_branch;
  wire T326;
  reg  ex_reg_branch;
  wire T327;
  wire id_branch;
  wire[31:0] T328;
  wire T329;
  wire ctrl_killx;
  wire T330;
  wire T331;
  reg  ex_reg_load_use;
  wire T332;
  wire id_load_use;
  wire T333;
  wire T334;
  wire replay_ex_structural;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  reg  mem_reg_sret;
  wire T340;
  reg  ex_reg_sret;
  wire T341;
  wire id_sret;
  wire[31:0] T342;
  wire ctrl_killm;
  wire T343;
  wire fpu_kill_mem;
  wire T344;
  wire killm_common;
  wire T345;
  reg  mem_reg_valid;
  wire T346;
  reg  ex_reg_valid;
  wire T347;
  wire T348;
  reg  mem_reg_xcpt;
  wire T349;
  wire ex_xcpt;
  wire T350;
  wire T351;
  reg  ex_reg_xcpt;
  wire T352;
  wire id_xcpt;
  wire id_syscall;
  wire[31:0] T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire id_csr_privileged;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire[1:0] T363;
  wire T364;
  wire T365;
  wire[1:0] T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire T372;
  wire T373;
  wire[1:0] T374;
  wire T375;
  wire T376;
  wire[1:0] T377;
  wire T378;
  wire T379;
  wire id_csr_invalid;
  wire T380;
  reg  T381;
  wire T383;
  wire id_int_val;
  wire T384;
  wire[31:0] T385;
  wire T386;
  wire T387;
  wire[31:0] T388;
  wire T389;
  wire T390;
  wire[31:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[31:0] T396;
  wire T397;
  wire T398;
  wire[31:0] T399;
  wire T400;
  wire T401;
  wire[31:0] T402;
  wire T403;
  wire T404;
  wire[31:0] T405;
  wire T406;
  wire T407;
  wire[31:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire[31:0] T412;
  wire T413;
  wire T414;
  wire[31:0] T415;
  wire T416;
  wire T417;
  wire[31:0] T418;
  wire T419;
  wire T420;
  wire[31:0] T421;
  wire T422;
  wire T423;
  wire[31:0] T424;
  wire T425;
  wire T426;
  wire[31:0] T427;
  wire T428;
  wire T429;
  wire[31:0] T430;
  wire T431;
  wire T432;
  wire[31:0] T433;
  wire T434;
  wire T435;
  wire[31:0] T436;
  wire T437;
  wire T438;
  wire[31:0] T439;
  wire T440;
  wire T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire[31:0] T445;
  wire T446;
  wire T447;
  wire T448;
  reg  ex_reg_xcpt_interrupt;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire dcache_kill_mem;
  wire T453;
  wire replay_wb;
  wire T454;
  wire T455;
  wire replay_wb_common;
  wire T456;
  reg  wb_reg_replay;
  wire T457;
  wire T458;
  wire replay_mem;
  wire T459;
  wire mem_xcpt;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  reg  mem_reg_xcpt_interrupt;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire wb_rocc_val;
  wire T472;
  wire T473;
  reg  wb_reg_flush_inst;
  wire T474;
  reg  mem_reg_flush_inst;
  wire T475;
  reg  ex_reg_flush_inst;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T483;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T484;
  wire T485;
  wire T486;
  reg  ex_reg_btb_hit;
  wire T487;
  reg [3:0] mem_reg_btb_resp_bht_index;
  wire[3:0] T488;
  reg [3:0] ex_reg_btb_resp_bht_index;
  wire[3:0] T489;
  reg [2:0] mem_reg_btb_resp_entry;
  wire[2:0] T490;
  reg [2:0] ex_reg_btb_resp_entry;
  wire[2:0] T491;
  reg [42:0] mem_reg_btb_resp_target;
  wire[42:0] T492;
  reg [42:0] ex_reg_btb_resp_target;
  wire[42:0] T493;
  reg  mem_reg_btb_resp_taken;
  wire T494;
  reg  ex_reg_btb_resp_taken;
  wire T495;
  reg  mem_reg_btb_hit;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  reg [63:0] wb_reg_cause;
  wire[63:0] T501;
  wire[63:0] mem_cause;
  wire[63:0] T667;
  wire[3:0] T502;
  wire[3:0] T503;
  wire[3:0] T504;
  reg [63:0] mem_reg_cause;
  wire[63:0] T505;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T506;
  wire[63:0] id_cause;
  wire[63:0] T668;
  wire[3:0] T507;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[3:0] T510;
  wire[3:0] T511;
  wire[3:0] T512;
  wire[63:0] id_interrupt_cause;
  wire[63:0] T513;
  wire[63:0] T514;
  wire[63:0] T515;
  wire[63:0] T516;
  wire[63:0] T517;
  wire[63:0] T518;
  wire T519;
  wire T520;
  reg  wb_reg_valid;
  wire T521;
  wire T522;
  wire[1:0] T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire[1:0] T533;
  wire[1:0] T534;
  wire[1:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire[2:0] T669;
  reg [1:0] wb_reg_csr;
  wire[1:0] T564;
  wire T565;
  wire[3:0] T566;
  wire[3:0] id_fn_alu;
  wire[2:0] T567;
  wire[1:0] T568;
  wire T569;
  wire T570;
  wire[31:0] T571;
  wire T572;
  wire T573;
  wire[31:0] T574;
  wire T575;
  wire[31:0] T576;
  wire T577;
  wire T578;
  wire[31:0] T579;
  wire T580;
  wire T581;
  wire[31:0] T582;
  wire T583;
  wire T584;
  wire[31:0] T585;
  wire T586;
  wire T587;
  wire[31:0] T588;
  wire T589;
  wire[31:0] T590;
  wire T591;
  wire T592;
  wire[31:0] T593;
  wire T594;
  wire T595;
  wire[31:0] T596;
  wire T597;
  wire T598;
  wire[31:0] T599;
  wire T600;
  wire[31:0] T601;
  wire T602;
  wire T603;
  wire[31:0] T604;
  wire T605;
  wire T606;
  wire T607;
  wire[31:0] T608;
  wire T609;
  wire id_fn_dw;
  wire T610;
  wire[31:0] T611;
  wire T612;
  wire[31:0] T613;
  wire[2:0] T614;
  wire[2:0] id_sel_imm;
  wire[1:0] T615;
  wire T616;
  wire T617;
  wire[31:0] T618;
  wire T619;
  wire[31:0] T620;
  wire T621;
  wire T622;
  wire[31:0] T623;
  wire T624;
  wire T625;
  wire[31:0] T626;
  wire T627;
  wire T628;
  wire[31:0] T629;
  wire[1:0] T630;
  wire[1:0] id_sel_alu1;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire[31:0] T635;
  wire T636;
  wire[31:0] T637;
  wire T638;
  wire T639;
  wire[31:0] T640;
  wire[2:0] T670;
  wire[1:0] T641;
  wire[1:0] id_sel_alu2;
  wire T642;
  wire T643;
  wire[31:0] T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire[31:0] T649;
  wire T650;
  wire[31:0] T651;
  wire T652;
  wire T653;
  wire[31:0] T654;
  wire T655;
  wire T656;
  wire T657;
  wire[31:0] T658;
  wire T659;
  wire T660;
  wire T661;
  wire[2:0] T671;
  wire[1:0] T662;
  wire[1:0] T663;
  wire[1:0] T664;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_xcpt = {1{$random}};
    wb_reg_sret = {1{$random}};
    mem_reg_replay = {1{$random}};
    mem_reg_replay_next = {1{$random}};
    ex_reg_replay_next = {1{$random}};
    id_reg_fence = {1{$random}};
    ex_reg_mem_val = {1{$random}};
    R105 = {1{$random}};
    wb_reg_rocc_val = {1{$random}};
    mem_reg_rocc_val = {1{$random}};
    ex_reg_rocc_val = {1{$random}};
    wb_reg_mem_val = {1{$random}};
    mem_reg_mem_val = {1{$random}};
    wb_reg_div_mul_val = {1{$random}};
    mem_reg_div_mul_val = {1{$random}};
    ex_reg_div_mul_val = {1{$random}};
    wb_reg_fp_val = {1{$random}};
    mem_reg_fp_val = {1{$random}};
    ex_reg_fp_val = {1{$random}};
    wb_reg_fp_wen = {1{$random}};
    mem_reg_fp_wen = {1{$random}};
    ex_reg_fp_wen = {1{$random}};
    wb_reg_wen = {1{$random}};
    mem_reg_wen = {1{$random}};
    ex_reg_wen = {1{$random}};
    mem_mem_cmd_bh = {1{$random}};
    ex_reg_mem_type = {1{$random}};
    ex_reg_mem_cmd = {1{$random}};
    mem_reg_csr = {1{$random}};
    ex_reg_csr = {1{$random}};
    ex_reg_jalr = {1{$random}};
    mem_reg_jal = {1{$random}};
    ex_reg_jal = {1{$random}};
    mem_reg_jalr = {1{$random}};
    mem_reg_branch = {1{$random}};
    ex_reg_branch = {1{$random}};
    ex_reg_load_use = {1{$random}};
    mem_reg_sret = {1{$random}};
    ex_reg_sret = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    wb_reg_replay = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    wb_reg_flush_inst = {1{$random}};
    mem_reg_flush_inst = {1{$random}};
    ex_reg_flush_inst = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_index = {1{$random}};
    ex_reg_btb_resp_bht_index = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_reg_valid = {1{$random}};
    wb_reg_csr = {1{$random}};
  end
`endif

  assign io_rocc_exception = T0;
  assign T0 = wb_reg_xcpt & io_dpath_status_er;
  assign T1 = mem_xcpt & T2;
  assign T2 = take_pc_wb ^ 1'h1;
  assign take_pc_wb = T3;
  assign T3 = T453 | wb_reg_sret;
  assign T4 = ctrl_killm ? 1'h0 : T5;
  assign T5 = mem_reg_sret & T6;
  assign T6 = mem_reg_replay ^ 1'h1;
  assign T7 = T339 & replay_ex;
  assign replay_ex = replay_ex_structural | replay_ex_other;
  assign replay_ex_other = T331 | mem_reg_replay_next;
  assign T8 = ctrl_killx ? 1'h0 : ex_reg_replay_next;
  assign T9 = ctrl_killd ? 1'h0 : T10;
  assign T10 = id_replay_next | id_csr_flush;
  assign id_csr_flush = T17 & T11;
  assign T11 = T12 ^ 1'h1;
  assign T12 = T15 | T13;
  assign T13 = T14 == 12'h0;
  assign T14 = id_csr_addr & 12'h88d;
  assign id_csr_addr = io_dpath_inst[5'h1f:5'h14];
  assign T15 = T16 == 12'h0;
  assign T16 = id_csr_addr & 12'h88e;
  assign T17 = id_csr_en & id_csr_wen;
  assign id_csr_wen = T26 | T18;
  assign T18 = T19 ^ 1'h1;
  assign T19 = T25 | T20;
  assign T20 = 2'h3 == id_csr;
  assign id_csr = {T23, T21};
  assign T21 = T22 == 32'h1050;
  assign T22 = io_dpath_inst & 32'h1050;
  assign T23 = T24 == 32'h2050;
  assign T24 = io_dpath_inst & 32'h2050;
  assign T25 = 2'h2 == id_csr;
  assign T26 = id_raddr1 != 5'h0;
  assign id_raddr1 = io_dpath_inst[5'h13:4'hf];
  assign id_csr_en = id_csr != 2'h0;
  assign id_replay_next = T27 == 32'h1008;
  assign T27 = io_dpath_inst & 32'h3058;
  assign ctrl_killd = T28;
  assign T28 = T59 | ctrl_draind;
  assign ctrl_draind = id_interrupt | ex_reg_replay_next;
  assign id_interrupt = io_dpath_status_ei & id_interrupt_unmasked;
  assign id_interrupt_unmasked = T32 | T29;
  assign T29 = T31 & T30;
  assign T30 = io_dpath_status_ip[3'h7:3'h7];
  assign T31 = io_dpath_status_im[3'h7:3'h7];
  assign T32 = T36 | T33;
  assign T33 = T35 & T34;
  assign T34 = io_dpath_status_ip[3'h6:3'h6];
  assign T35 = io_dpath_status_im[3'h6:3'h6];
  assign T36 = T40 | T37;
  assign T37 = T39 & T38;
  assign T38 = io_dpath_status_ip[3'h5:3'h5];
  assign T39 = io_dpath_status_im[3'h5:3'h5];
  assign T40 = T44 | T41;
  assign T41 = T43 & T42;
  assign T42 = io_dpath_status_ip[3'h4:3'h4];
  assign T43 = io_dpath_status_im[3'h4:3'h4];
  assign T44 = T48 | T45;
  assign T45 = T47 & T46;
  assign T46 = io_dpath_status_ip[2'h3:2'h3];
  assign T47 = io_dpath_status_im[2'h3:2'h3];
  assign T48 = T52 | T49;
  assign T49 = T51 & T50;
  assign T50 = io_dpath_status_ip[2'h2:2'h2];
  assign T51 = io_dpath_status_im[2'h2:2'h2];
  assign T52 = T56 | T53;
  assign T53 = T55 & T54;
  assign T54 = io_dpath_status_ip[1'h1:1'h1];
  assign T55 = io_dpath_status_im[1'h1:1'h1];
  assign T56 = T58 & T57;
  assign T57 = io_dpath_status_ip[1'h0:1'h0];
  assign T58 = io_dpath_status_im[1'h0:1'h0];
  assign T59 = T320 | ctrl_stalld;
  assign ctrl_stalld = T90 | id_do_fence;
  assign id_do_fence = id_mem_busy & T60;
  assign T60 = T61 | id_csr_flush;
  assign T61 = T84 | T62;
  assign T62 = id_reg_fence & id_mem_val;
  assign id_mem_val = T65 | T63;
  assign T63 = T64 == 32'h1000202f;
  assign T64 = io_dpath_inst & 32'hf9f0607f;
  assign T65 = T68 | T66;
  assign T66 = T67 == 32'h800202f;
  assign T67 = io_dpath_inst & 32'he800607f;
  assign T68 = T71 | T69;
  assign T69 = T70 == 32'h202f;
  assign T70 = io_dpath_inst & 32'h1800607f;
  assign T71 = T74 | T72;
  assign T72 = T73 == 32'h3;
  assign T73 = io_dpath_inst & 32'h107f;
  assign T74 = T77 | T75;
  assign T75 = T76 == 32'h3;
  assign T76 = io_dpath_inst & 32'h207f;
  assign T77 = T78 == 32'h3;
  assign T78 = io_dpath_inst & 32'h405f;
  assign T665 = reset ? 1'h0 : T79;
  assign T79 = id_fence_next | T80;
  assign T80 = id_reg_fence & id_mem_busy;
  assign id_fence_next = id_fence | T81;
  assign T81 = id_amo & id_amo_rl;
  assign id_amo_rl = io_dpath_inst[5'h19:5'h19];
  assign id_amo = T82 == 32'h2008;
  assign T82 = io_dpath_inst & 32'h6048;
  assign id_fence = T83 == 32'h8;
  assign T83 = io_dpath_inst & 32'h3058;
  assign T84 = T86 | id_fence_i;
  assign id_fence_i = T85 == 32'h100f;
  assign T85 = io_dpath_inst & 32'h707f;
  assign T86 = id_amo & id_amo_aq;
  assign id_amo_aq = io_dpath_inst[5'h1a:5'h1a];
  assign id_mem_busy = T89 | ex_reg_mem_val;
  assign T87 = ctrl_killd ? 1'h0 : T88;
  assign T88 = id_mem_val;
  assign T89 = io_dmem_ordered ^ 1'h1;
  assign T90 = T93 | T91;
  assign T91 = id_mem_val & T92;
  assign T92 = io_dmem_req_ready ^ 1'h1;
  assign T93 = T183 | id_sboard_hazard;
  assign id_sboard_hazard = T146 | T94;
  assign T94 = id_wen_not0 & T95;
  assign T95 = T100 & T96;
  assign T96 = T97 - 1'h1;
  assign T97 = 1'h1 << T98;
  assign T98 = T99 + 5'h1;
  assign T99 = id_waddr - id_waddr;
  assign id_waddr = io_dpath_inst[4'hb:3'h7];
  assign T100 = T101 >> id_waddr;
  assign T101 = R105 & T102;
  assign T102 = ~ T103;
  assign T103 = io_dpath_ll_wen ? T104 : 32'h0;
  assign T104 = 1'h1 << io_dpath_ll_waddr;
  assign T666 = reset ? 32'h0 : T106;
  assign T106 = T126 ? T108 : T107;
  assign T107 = io_dpath_ll_wen ? T101 : R105;
  assign T108 = T101 | T109;
  assign T109 = T111 ? T110 : 32'h0;
  assign T110 = 1'h1 << io_dpath_wb_waddr;
  assign T111 = wb_set_sboard & io_dpath_wb_wen;
  assign wb_set_sboard = T116 | wb_reg_rocc_val;
  assign T112 = ctrl_killm ? 1'h0 : mem_reg_rocc_val;
  assign T113 = ctrl_killx ? 1'h0 : ex_reg_rocc_val;
  assign T114 = ctrl_killd ? 1'h0 : T115;
  assign T115 = 1'h0;
  assign T116 = wb_reg_div_mul_val | wb_dcache_miss;
  assign wb_dcache_miss = wb_reg_mem_val & T117;
  assign T117 = io_dmem_resp_valid ^ 1'h1;
  assign T118 = ctrl_killm ? 1'h0 : mem_reg_mem_val;
  assign T119 = ctrl_killx ? 1'h0 : ex_reg_mem_val;
  assign T120 = ctrl_killm ? 1'h0 : mem_reg_div_mul_val;
  assign T121 = ex_reg_div_mul_val & io_dpath_div_mul_rdy;
  assign T122 = ctrl_killd ? 1'h0 : T123;
  assign T123 = id_mul_val | id_div_val;
  assign id_div_val = T124 == 32'h2004020;
  assign T124 = io_dpath_inst & 32'h2004064;
  assign id_mul_val = T125 == 32'h2000030;
  assign T125 = io_dpath_inst & 32'h2004074;
  assign T126 = io_dpath_ll_wen | T111;
  assign id_wen_not0 = id_wen & T127;
  assign T127 = id_waddr != 5'h0;
  assign id_wen = T130 | T128;
  assign T128 = T129 == 32'h0;
  assign T129 = io_dpath_inst & 32'h28;
  assign T130 = T133 | T131;
  assign T131 = T132 == 32'h2010;
  assign T132 = io_dpath_inst & 32'h2010;
  assign T133 = T136 | T134;
  assign T134 = T135 == 32'h2008;
  assign T135 = io_dpath_inst & 32'h2008;
  assign T136 = T139 | T137;
  assign T137 = T138 == 32'h1010;
  assign T138 = io_dpath_inst & 32'h1010;
  assign T139 = T141 | id_jal;
  assign id_jal = T140 == 32'h48;
  assign T140 = io_dpath_inst & 32'h48;
  assign T141 = T144 | T142;
  assign T142 = T143 == 32'h10;
  assign T143 = io_dpath_inst & 32'h50;
  assign T144 = T145 == 32'h4;
  assign T145 = io_dpath_inst & 32'hc;
  assign T146 = T162 | T147;
  assign T147 = id_renx2_not0 & T148;
  assign T148 = T153 & T149;
  assign T149 = T150 - 1'h1;
  assign T150 = 1'h1 << T151;
  assign T151 = T152 + 5'h1;
  assign T152 = id_raddr2 - id_raddr2;
  assign id_raddr2 = io_dpath_inst[5'h18:5'h14];
  assign T153 = T101 >> id_raddr2;
  assign id_renx2_not0 = id_renx2 & T154;
  assign T154 = id_raddr2 != 5'h0;
  assign id_renx2 = T157 | T155;
  assign T155 = T156 == 32'h20;
  assign T156 = io_dpath_inst & 32'h34;
  assign T157 = T160 | T158;
  assign T158 = T159 == 32'h20;
  assign T159 = io_dpath_inst & 32'h64;
  assign T160 = T161 == 32'h20;
  assign T161 = io_dpath_inst & 32'h70;
  assign T162 = id_renx1_not0 & T163;
  assign T163 = T168 & T164;
  assign T164 = T165 - 1'h1;
  assign T165 = 1'h1 << T166;
  assign T166 = T167 + 5'h1;
  assign T167 = id_raddr1 - id_raddr1;
  assign T168 = T101 >> id_raddr1;
  assign id_renx1_not0 = id_renx1 & T169;
  assign T169 = id_raddr1 != 5'h0;
  assign id_renx1 = T172 | T170;
  assign T170 = T171 == 32'h2000;
  assign T171 = io_dpath_inst & 32'h2050;
  assign T172 = T175 | T173;
  assign T173 = T174 == 32'h2000;
  assign T174 = io_dpath_inst & 32'h6004;
  assign T175 = T178 | T176;
  assign T176 = T177 == 32'h1000;
  assign T177 = io_dpath_inst & 32'h5004;
  assign T178 = T181 | T179;
  assign T179 = T180 == 32'h0;
  assign T180 = io_dpath_inst & 32'h18;
  assign T181 = T182 == 32'h0;
  assign T182 = io_dpath_inst & 32'h44;
  assign T183 = T215 | id_wb_hazard;
  assign id_wb_hazard = T203 | T184;
  assign T184 = fp_data_hazard_wb & T185;
  assign T185 = wb_dcache_miss | wb_reg_fp_val;
  assign T186 = ctrl_killm ? 1'h0 : mem_reg_fp_val;
  assign T187 = ctrl_killx ? 1'h0 : ex_reg_fp_val;
  assign T188 = ctrl_killd ? 1'h0 : 1'h0;
  assign fp_data_hazard_wb = wb_reg_fp_wen & T189;
  assign T189 = T192 | T190;
  assign T190 = io_fpu_dec_wen & T191;
  assign T191 = id_waddr == io_dpath_wb_waddr;
  assign T192 = T195 | T193;
  assign T193 = io_fpu_dec_ren3 & T194;
  assign T194 = id_raddr3 == io_dpath_wb_waddr;
  assign id_raddr3 = io_dpath_inst[5'h1f:5'h1b];
  assign T195 = T198 | T196;
  assign T196 = io_fpu_dec_ren2 & T197;
  assign T197 = id_raddr2 == io_dpath_wb_waddr;
  assign T198 = io_fpu_dec_ren1 & T199;
  assign T199 = id_raddr1 == io_dpath_wb_waddr;
  assign T200 = ctrl_killm ? 1'h0 : mem_reg_fp_wen;
  assign T201 = ctrl_killx ? 1'h0 : ex_reg_fp_wen;
  assign T202 = ctrl_killd ? 1'h0 : 1'h0;
  assign T203 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_reg_wen & T204;
  assign T204 = T207 | T205;
  assign T205 = id_wen_not0 & T206;
  assign T206 = id_waddr == io_dpath_wb_waddr;
  assign T207 = T210 | T208;
  assign T208 = id_renx2_not0 & T209;
  assign T209 = id_raddr2 == io_dpath_wb_waddr;
  assign T210 = id_renx1_not0 & T211;
  assign T211 = id_raddr1 == io_dpath_wb_waddr;
  assign T212 = ctrl_killm ? 1'h0 : mem_reg_wen;
  assign T213 = ctrl_killx ? 1'h0 : ex_reg_wen;
  assign T214 = ctrl_killd ? 1'h0 : id_wen;
  assign T215 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = T228 | T216;
  assign T216 = fp_data_hazard_mem & mem_reg_fp_val;
  assign fp_data_hazard_mem = mem_reg_fp_wen & T217;
  assign T217 = T220 | T218;
  assign T218 = io_fpu_dec_wen & T219;
  assign T219 = id_waddr == io_dpath_mem_waddr;
  assign T220 = T223 | T221;
  assign T221 = io_fpu_dec_ren3 & T222;
  assign T222 = id_raddr3 == io_dpath_mem_waddr;
  assign T223 = T226 | T224;
  assign T224 = io_fpu_dec_ren2 & T225;
  assign T225 = id_raddr2 == io_dpath_mem_waddr;
  assign T226 = io_fpu_dec_ren1 & T227;
  assign T227 = id_raddr1 == io_dpath_mem_waddr;
  assign T228 = data_hazard_mem & T229;
  assign T229 = T230 | mem_reg_rocc_val;
  assign T230 = T231 | mem_reg_fp_val;
  assign T231 = T232 | mem_reg_div_mul_val;
  assign T232 = T279 | T233;
  assign T233 = mem_reg_mem_val & mem_mem_cmd_bh;
  assign T234 = T278 ? ex_slow_bypass : mem_mem_cmd_bh;
  assign ex_slow_bypass = T252 | T235;
  assign T235 = T247 | T236;
  assign T236 = 3'h5 == ex_reg_mem_type;
  assign T237 = T246 ? T238 : ex_reg_mem_type;
  assign T238 = id_mem_type;
  assign id_mem_type = {T244, T239};
  assign T239 = {T242, T240};
  assign T240 = T241 == 32'h1000;
  assign T241 = io_dpath_inst & 32'h1000;
  assign T242 = T243 == 32'h2000;
  assign T243 = io_dpath_inst & 32'h2000;
  assign T244 = T245 == 32'h4000;
  assign T245 = io_dpath_inst & 32'h4000;
  assign T246 = ctrl_killd ^ 1'h1;
  assign T247 = T249 | T248;
  assign T248 = 3'h1 == ex_reg_mem_type;
  assign T249 = T251 | T250;
  assign T250 = 3'h4 == ex_reg_mem_type;
  assign T251 = 3'h0 == ex_reg_mem_type;
  assign T252 = ex_reg_mem_cmd == 5'h7;
  assign T253 = T246 ? id_mem_cmd : ex_reg_mem_cmd;
  assign id_mem_cmd = {1'h0, T254};
  assign T254 = {T276, T255};
  assign T255 = {T270, T256};
  assign T256 = {T265, T257};
  assign T257 = T260 | T258;
  assign T258 = T259 == 32'h20000020;
  assign T259 = io_dpath_inst & 32'h20000020;
  assign T260 = T263 | T261;
  assign T261 = T262 == 32'h18000020;
  assign T262 = io_dpath_inst & 32'h18000020;
  assign T263 = T264 == 32'h20;
  assign T264 = io_dpath_inst & 32'h28;
  assign T265 = T268 | T266;
  assign T266 = T267 == 32'h40000008;
  assign T267 = io_dpath_inst & 32'h40000008;
  assign T268 = T269 == 32'h10000008;
  assign T269 = io_dpath_inst & 32'h10000008;
  assign T270 = T273 | T271;
  assign T271 = T272 == 32'h80000008;
  assign T272 = io_dpath_inst & 32'h80000008;
  assign T273 = T274 | T268;
  assign T274 = T275 == 32'h8000008;
  assign T275 = io_dpath_inst & 32'h8000008;
  assign T276 = T277 == 32'h8;
  assign T277 = io_dpath_inst & 32'h18000008;
  assign T278 = ctrl_killx ^ 1'h1;
  assign T279 = mem_reg_csr != 2'h0;
  assign T280 = ctrl_killx ? 2'h0 : ex_reg_csr;
  assign T281 = ctrl_killd ? 2'h0 : id_csr;
  assign data_hazard_mem = mem_reg_wen & T282;
  assign T282 = T285 | T283;
  assign T283 = id_wen_not0 & T284;
  assign T284 = id_waddr == io_dpath_mem_waddr;
  assign T285 = T288 | T286;
  assign T286 = id_renx2_not0 & T287;
  assign T287 = id_raddr2 == io_dpath_mem_waddr;
  assign T288 = id_renx1_not0 & T289;
  assign T289 = id_raddr1 == io_dpath_mem_waddr;
  assign id_ex_hazard = T303 | T290;
  assign T290 = fp_data_hazard_ex & T291;
  assign T291 = ex_reg_mem_val | ex_reg_fp_val;
  assign fp_data_hazard_ex = ex_reg_fp_wen & T292;
  assign T292 = T295 | T293;
  assign T293 = io_fpu_dec_wen & T294;
  assign T294 = id_waddr == io_dpath_ex_waddr;
  assign T295 = T298 | T296;
  assign T296 = io_fpu_dec_ren3 & T297;
  assign T297 = id_raddr3 == io_dpath_ex_waddr;
  assign T298 = T301 | T299;
  assign T299 = io_fpu_dec_ren2 & T300;
  assign T300 = id_raddr2 == io_dpath_ex_waddr;
  assign T301 = io_fpu_dec_ren1 & T302;
  assign T302 = id_raddr1 == io_dpath_ex_waddr;
  assign T303 = data_hazard_ex & T304;
  assign T304 = T305 | ex_reg_rocc_val;
  assign T305 = T306 | ex_reg_fp_val;
  assign T306 = T307 | ex_reg_div_mul_val;
  assign T307 = T308 | ex_reg_mem_val;
  assign T308 = T311 | ex_reg_jalr;
  assign T309 = ctrl_killd ? 1'h0 : id_jalr;
  assign id_jalr = T310 == 32'h4;
  assign T310 = io_dpath_inst & 32'h1c;
  assign T311 = ex_reg_csr != 2'h0;
  assign data_hazard_ex = ex_reg_wen & T312;
  assign T312 = T315 | T313;
  assign T313 = id_wen_not0 & T314;
  assign T314 = id_waddr == io_dpath_ex_waddr;
  assign T315 = T318 | T316;
  assign T316 = id_renx2_not0 & T317;
  assign T317 = id_raddr2 == io_dpath_ex_waddr;
  assign T318 = id_renx1_not0 & T319;
  assign T319 = id_raddr1 == io_dpath_ex_waddr;
  assign T320 = T329 | take_pc;
  assign take_pc = take_pc_wb | take_pc_mem;
  assign take_pc_mem = io_dpath_mem_misprediction & T321;
  assign T321 = T324 | mem_reg_jal;
  assign T322 = ctrl_killx ? 1'h0 : ex_reg_jal;
  assign T323 = ctrl_killd ? 1'h0 : id_jal;
  assign T324 = mem_reg_branch | mem_reg_jalr;
  assign T325 = ctrl_killx ? 1'h0 : ex_reg_jalr;
  assign T326 = ctrl_killx ? 1'h0 : ex_reg_branch;
  assign T327 = ctrl_killd ? 1'h0 : id_branch;
  assign id_branch = T328 == 32'h40;
  assign T328 = io_dpath_inst & 32'h54;
  assign T329 = io_imem_resp_valid ^ 1'h1;
  assign ctrl_killx = T330;
  assign T330 = take_pc | replay_ex;
  assign T331 = wb_dcache_miss & ex_reg_load_use;
  assign T332 = ctrl_killd ? 1'h0 : id_load_use;
  assign id_load_use = T333;
  assign T333 = mem_reg_mem_val & T334;
  assign T334 = data_hazard_mem | fp_data_hazard_mem;
  assign replay_ex_structural = T337 | T335;
  assign T335 = ex_reg_div_mul_val & T336;
  assign T336 = io_dpath_div_mul_rdy ^ 1'h1;
  assign T337 = ex_reg_mem_val & T338;
  assign T338 = io_dmem_req_ready ^ 1'h1;
  assign T339 = take_pc ^ 1'h1;
  assign T340 = ctrl_killx ? 1'h0 : ex_reg_sret;
  assign T341 = ctrl_killd ? 1'h0 : id_sret;
  assign id_sret = T342 == 32'h80000050;
  assign T342 = io_dpath_inst & 32'h80003050;
  assign ctrl_killm = T343;
  assign T343 = T344 | fpu_kill_mem;
  assign fpu_kill_mem = mem_reg_fp_val & io_fpu_nack_mem;
  assign T344 = killm_common | mem_xcpt;
  assign killm_common = T348 | T345;
  assign T345 = mem_reg_valid ^ 1'h1;
  assign T346 = ctrl_killx ? 1'h0 : ex_reg_valid;
  assign T347 = ctrl_killd ? 1'h0 : 1'h1;
  assign T348 = T452 | mem_reg_xcpt;
  assign T349 = ctrl_killx ? 1'h0 : ex_xcpt;
  assign ex_xcpt = T351 | T350;
  assign T350 = ex_reg_fp_val & io_fpu_illegal_rm;
  assign T351 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T352 = ctrl_killd ? 1'h0 : id_xcpt;
  assign id_xcpt = T354 | id_syscall;
  assign id_syscall = T353 == 32'h50;
  assign T353 = io_dpath_inst & 32'h80003050;
  assign T354 = T357 | T355;
  assign T355 = id_sret & T356;
  assign T356 = io_dpath_status_s ^ 1'h1;
  assign T357 = T378 | id_csr_privileged;
  assign id_csr_privileged = id_csr_en & T358;
  assign T358 = T364 | T359;
  assign T359 = T360 & id_csr_wen;
  assign T360 = T362 & T361;
  assign T361 = io_dpath_status_s ^ 1'h1;
  assign T362 = T363 == 2'h1;
  assign T363 = id_csr_addr[4'h9:4'h8];
  assign T364 = T367 | T365;
  assign T365 = 2'h2 <= T366;
  assign T366 = id_csr_addr[4'h9:4'h8];
  assign T367 = T372 | T368;
  assign T368 = T370 & T369;
  assign T369 = io_dpath_status_s ^ 1'h1;
  assign T370 = T371 == 2'h1;
  assign T371 = id_csr_addr[4'hb:4'ha];
  assign T372 = T375 | T373;
  assign T373 = T374 == 2'h2;
  assign T374 = id_csr_addr[4'hb:4'ha];
  assign T375 = T376 & id_csr_wen;
  assign T376 = T377 == 2'h3;
  assign T377 = id_csr_addr[4'hb:4'ha];
  assign T378 = T447 | T379;
  assign T379 = T383 | id_csr_invalid;
  assign id_csr_invalid = id_csr_en & T380;
  assign T380 = T381 ^ 1'h1;
  always @(*) case (id_csr_addr)
    0: T381 = 1'h0;
    1: T381 = 1'h0;
    2: T381 = 1'h0;
    3: T381 = 1'h0;
    4: T381 = 1'h0;
    5: T381 = 1'h0;
    6: T381 = 1'h0;
    7: T381 = 1'h0;
    8: T381 = 1'h0;
    9: T381 = 1'h0;
    10: T381 = 1'h0;
    11: T381 = 1'h0;
    12: T381 = 1'h0;
    13: T381 = 1'h0;
    14: T381 = 1'h0;
    15: T381 = 1'h0;
    16: T381 = 1'h0;
    17: T381 = 1'h0;
    18: T381 = 1'h0;
    19: T381 = 1'h0;
    20: T381 = 1'h0;
    21: T381 = 1'h0;
    22: T381 = 1'h0;
    23: T381 = 1'h0;
    24: T381 = 1'h0;
    25: T381 = 1'h0;
    26: T381 = 1'h0;
    27: T381 = 1'h0;
    28: T381 = 1'h0;
    29: T381 = 1'h0;
    30: T381 = 1'h0;
    31: T381 = 1'h0;
    32: T381 = 1'h0;
    33: T381 = 1'h0;
    34: T381 = 1'h0;
    35: T381 = 1'h0;
    36: T381 = 1'h0;
    37: T381 = 1'h0;
    38: T381 = 1'h0;
    39: T381 = 1'h0;
    40: T381 = 1'h0;
    41: T381 = 1'h0;
    42: T381 = 1'h0;
    43: T381 = 1'h0;
    44: T381 = 1'h0;
    45: T381 = 1'h0;
    46: T381 = 1'h0;
    47: T381 = 1'h0;
    48: T381 = 1'h0;
    49: T381 = 1'h0;
    50: T381 = 1'h0;
    51: T381 = 1'h0;
    52: T381 = 1'h0;
    53: T381 = 1'h0;
    54: T381 = 1'h0;
    55: T381 = 1'h0;
    56: T381 = 1'h0;
    57: T381 = 1'h0;
    58: T381 = 1'h0;
    59: T381 = 1'h0;
    60: T381 = 1'h0;
    61: T381 = 1'h0;
    62: T381 = 1'h0;
    63: T381 = 1'h0;
    64: T381 = 1'h0;
    65: T381 = 1'h0;
    66: T381 = 1'h0;
    67: T381 = 1'h0;
    68: T381 = 1'h0;
    69: T381 = 1'h0;
    70: T381 = 1'h0;
    71: T381 = 1'h0;
    72: T381 = 1'h0;
    73: T381 = 1'h0;
    74: T381 = 1'h0;
    75: T381 = 1'h0;
    76: T381 = 1'h0;
    77: T381 = 1'h0;
    78: T381 = 1'h0;
    79: T381 = 1'h0;
    80: T381 = 1'h0;
    81: T381 = 1'h0;
    82: T381 = 1'h0;
    83: T381 = 1'h0;
    84: T381 = 1'h0;
    85: T381 = 1'h0;
    86: T381 = 1'h0;
    87: T381 = 1'h0;
    88: T381 = 1'h0;
    89: T381 = 1'h0;
    90: T381 = 1'h0;
    91: T381 = 1'h0;
    92: T381 = 1'h0;
    93: T381 = 1'h0;
    94: T381 = 1'h0;
    95: T381 = 1'h0;
    96: T381 = 1'h0;
    97: T381 = 1'h0;
    98: T381 = 1'h0;
    99: T381 = 1'h0;
    100: T381 = 1'h0;
    101: T381 = 1'h0;
    102: T381 = 1'h0;
    103: T381 = 1'h0;
    104: T381 = 1'h0;
    105: T381 = 1'h0;
    106: T381 = 1'h0;
    107: T381 = 1'h0;
    108: T381 = 1'h0;
    109: T381 = 1'h0;
    110: T381 = 1'h0;
    111: T381 = 1'h0;
    112: T381 = 1'h0;
    113: T381 = 1'h0;
    114: T381 = 1'h0;
    115: T381 = 1'h0;
    116: T381 = 1'h0;
    117: T381 = 1'h0;
    118: T381 = 1'h0;
    119: T381 = 1'h0;
    120: T381 = 1'h0;
    121: T381 = 1'h0;
    122: T381 = 1'h0;
    123: T381 = 1'h0;
    124: T381 = 1'h0;
    125: T381 = 1'h0;
    126: T381 = 1'h0;
    127: T381 = 1'h0;
    128: T381 = 1'h0;
    129: T381 = 1'h0;
    130: T381 = 1'h0;
    131: T381 = 1'h0;
    132: T381 = 1'h0;
    133: T381 = 1'h0;
    134: T381 = 1'h0;
    135: T381 = 1'h0;
    136: T381 = 1'h0;
    137: T381 = 1'h0;
    138: T381 = 1'h0;
    139: T381 = 1'h0;
    140: T381 = 1'h0;
    141: T381 = 1'h0;
    142: T381 = 1'h0;
    143: T381 = 1'h0;
    144: T381 = 1'h0;
    145: T381 = 1'h0;
    146: T381 = 1'h0;
    147: T381 = 1'h0;
    148: T381 = 1'h0;
    149: T381 = 1'h0;
    150: T381 = 1'h0;
    151: T381 = 1'h0;
    152: T381 = 1'h0;
    153: T381 = 1'h0;
    154: T381 = 1'h0;
    155: T381 = 1'h0;
    156: T381 = 1'h0;
    157: T381 = 1'h0;
    158: T381 = 1'h0;
    159: T381 = 1'h0;
    160: T381 = 1'h0;
    161: T381 = 1'h0;
    162: T381 = 1'h0;
    163: T381 = 1'h0;
    164: T381 = 1'h0;
    165: T381 = 1'h0;
    166: T381 = 1'h0;
    167: T381 = 1'h0;
    168: T381 = 1'h0;
    169: T381 = 1'h0;
    170: T381 = 1'h0;
    171: T381 = 1'h0;
    172: T381 = 1'h0;
    173: T381 = 1'h0;
    174: T381 = 1'h0;
    175: T381 = 1'h0;
    176: T381 = 1'h0;
    177: T381 = 1'h0;
    178: T381 = 1'h0;
    179: T381 = 1'h0;
    180: T381 = 1'h0;
    181: T381 = 1'h0;
    182: T381 = 1'h0;
    183: T381 = 1'h0;
    184: T381 = 1'h0;
    185: T381 = 1'h0;
    186: T381 = 1'h0;
    187: T381 = 1'h0;
    188: T381 = 1'h0;
    189: T381 = 1'h0;
    190: T381 = 1'h0;
    191: T381 = 1'h0;
    192: T381 = 1'h1;
    193: T381 = 1'h0;
    194: T381 = 1'h0;
    195: T381 = 1'h0;
    196: T381 = 1'h0;
    197: T381 = 1'h0;
    198: T381 = 1'h0;
    199: T381 = 1'h0;
    200: T381 = 1'h0;
    201: T381 = 1'h0;
    202: T381 = 1'h0;
    203: T381 = 1'h0;
    204: T381 = 1'h0;
    205: T381 = 1'h0;
    206: T381 = 1'h0;
    207: T381 = 1'h0;
    208: T381 = 1'h0;
    209: T381 = 1'h0;
    210: T381 = 1'h0;
    211: T381 = 1'h0;
    212: T381 = 1'h0;
    213: T381 = 1'h0;
    214: T381 = 1'h0;
    215: T381 = 1'h0;
    216: T381 = 1'h0;
    217: T381 = 1'h0;
    218: T381 = 1'h0;
    219: T381 = 1'h0;
    220: T381 = 1'h0;
    221: T381 = 1'h0;
    222: T381 = 1'h0;
    223: T381 = 1'h0;
    224: T381 = 1'h0;
    225: T381 = 1'h0;
    226: T381 = 1'h0;
    227: T381 = 1'h0;
    228: T381 = 1'h0;
    229: T381 = 1'h0;
    230: T381 = 1'h0;
    231: T381 = 1'h0;
    232: T381 = 1'h0;
    233: T381 = 1'h0;
    234: T381 = 1'h0;
    235: T381 = 1'h0;
    236: T381 = 1'h0;
    237: T381 = 1'h0;
    238: T381 = 1'h0;
    239: T381 = 1'h0;
    240: T381 = 1'h0;
    241: T381 = 1'h0;
    242: T381 = 1'h0;
    243: T381 = 1'h0;
    244: T381 = 1'h0;
    245: T381 = 1'h0;
    246: T381 = 1'h0;
    247: T381 = 1'h0;
    248: T381 = 1'h0;
    249: T381 = 1'h0;
    250: T381 = 1'h0;
    251: T381 = 1'h0;
    252: T381 = 1'h0;
    253: T381 = 1'h0;
    254: T381 = 1'h0;
    255: T381 = 1'h0;
    256: T381 = 1'h0;
    257: T381 = 1'h0;
    258: T381 = 1'h0;
    259: T381 = 1'h0;
    260: T381 = 1'h0;
    261: T381 = 1'h0;
    262: T381 = 1'h0;
    263: T381 = 1'h0;
    264: T381 = 1'h0;
    265: T381 = 1'h0;
    266: T381 = 1'h0;
    267: T381 = 1'h0;
    268: T381 = 1'h0;
    269: T381 = 1'h0;
    270: T381 = 1'h0;
    271: T381 = 1'h0;
    272: T381 = 1'h0;
    273: T381 = 1'h0;
    274: T381 = 1'h0;
    275: T381 = 1'h0;
    276: T381 = 1'h0;
    277: T381 = 1'h0;
    278: T381 = 1'h0;
    279: T381 = 1'h0;
    280: T381 = 1'h0;
    281: T381 = 1'h0;
    282: T381 = 1'h0;
    283: T381 = 1'h0;
    284: T381 = 1'h0;
    285: T381 = 1'h0;
    286: T381 = 1'h0;
    287: T381 = 1'h0;
    288: T381 = 1'h0;
    289: T381 = 1'h0;
    290: T381 = 1'h0;
    291: T381 = 1'h0;
    292: T381 = 1'h0;
    293: T381 = 1'h0;
    294: T381 = 1'h0;
    295: T381 = 1'h0;
    296: T381 = 1'h0;
    297: T381 = 1'h0;
    298: T381 = 1'h0;
    299: T381 = 1'h0;
    300: T381 = 1'h0;
    301: T381 = 1'h0;
    302: T381 = 1'h0;
    303: T381 = 1'h0;
    304: T381 = 1'h0;
    305: T381 = 1'h0;
    306: T381 = 1'h0;
    307: T381 = 1'h0;
    308: T381 = 1'h0;
    309: T381 = 1'h0;
    310: T381 = 1'h0;
    311: T381 = 1'h0;
    312: T381 = 1'h0;
    313: T381 = 1'h0;
    314: T381 = 1'h0;
    315: T381 = 1'h0;
    316: T381 = 1'h0;
    317: T381 = 1'h0;
    318: T381 = 1'h0;
    319: T381 = 1'h0;
    320: T381 = 1'h0;
    321: T381 = 1'h0;
    322: T381 = 1'h0;
    323: T381 = 1'h0;
    324: T381 = 1'h0;
    325: T381 = 1'h0;
    326: T381 = 1'h0;
    327: T381 = 1'h0;
    328: T381 = 1'h0;
    329: T381 = 1'h0;
    330: T381 = 1'h0;
    331: T381 = 1'h0;
    332: T381 = 1'h0;
    333: T381 = 1'h0;
    334: T381 = 1'h0;
    335: T381 = 1'h0;
    336: T381 = 1'h0;
    337: T381 = 1'h0;
    338: T381 = 1'h0;
    339: T381 = 1'h0;
    340: T381 = 1'h0;
    341: T381 = 1'h0;
    342: T381 = 1'h0;
    343: T381 = 1'h0;
    344: T381 = 1'h0;
    345: T381 = 1'h0;
    346: T381 = 1'h0;
    347: T381 = 1'h0;
    348: T381 = 1'h0;
    349: T381 = 1'h0;
    350: T381 = 1'h0;
    351: T381 = 1'h0;
    352: T381 = 1'h0;
    353: T381 = 1'h0;
    354: T381 = 1'h0;
    355: T381 = 1'h0;
    356: T381 = 1'h0;
    357: T381 = 1'h0;
    358: T381 = 1'h0;
    359: T381 = 1'h0;
    360: T381 = 1'h0;
    361: T381 = 1'h0;
    362: T381 = 1'h0;
    363: T381 = 1'h0;
    364: T381 = 1'h0;
    365: T381 = 1'h0;
    366: T381 = 1'h0;
    367: T381 = 1'h0;
    368: T381 = 1'h0;
    369: T381 = 1'h0;
    370: T381 = 1'h0;
    371: T381 = 1'h0;
    372: T381 = 1'h0;
    373: T381 = 1'h0;
    374: T381 = 1'h0;
    375: T381 = 1'h0;
    376: T381 = 1'h0;
    377: T381 = 1'h0;
    378: T381 = 1'h0;
    379: T381 = 1'h0;
    380: T381 = 1'h0;
    381: T381 = 1'h0;
    382: T381 = 1'h0;
    383: T381 = 1'h0;
    384: T381 = 1'h0;
    385: T381 = 1'h0;
    386: T381 = 1'h0;
    387: T381 = 1'h0;
    388: T381 = 1'h0;
    389: T381 = 1'h0;
    390: T381 = 1'h0;
    391: T381 = 1'h0;
    392: T381 = 1'h0;
    393: T381 = 1'h0;
    394: T381 = 1'h0;
    395: T381 = 1'h0;
    396: T381 = 1'h0;
    397: T381 = 1'h0;
    398: T381 = 1'h0;
    399: T381 = 1'h0;
    400: T381 = 1'h0;
    401: T381 = 1'h0;
    402: T381 = 1'h0;
    403: T381 = 1'h0;
    404: T381 = 1'h0;
    405: T381 = 1'h0;
    406: T381 = 1'h0;
    407: T381 = 1'h0;
    408: T381 = 1'h0;
    409: T381 = 1'h0;
    410: T381 = 1'h0;
    411: T381 = 1'h0;
    412: T381 = 1'h0;
    413: T381 = 1'h0;
    414: T381 = 1'h0;
    415: T381 = 1'h0;
    416: T381 = 1'h0;
    417: T381 = 1'h0;
    418: T381 = 1'h0;
    419: T381 = 1'h0;
    420: T381 = 1'h0;
    421: T381 = 1'h0;
    422: T381 = 1'h0;
    423: T381 = 1'h0;
    424: T381 = 1'h0;
    425: T381 = 1'h0;
    426: T381 = 1'h0;
    427: T381 = 1'h0;
    428: T381 = 1'h0;
    429: T381 = 1'h0;
    430: T381 = 1'h0;
    431: T381 = 1'h0;
    432: T381 = 1'h0;
    433: T381 = 1'h0;
    434: T381 = 1'h0;
    435: T381 = 1'h0;
    436: T381 = 1'h0;
    437: T381 = 1'h0;
    438: T381 = 1'h0;
    439: T381 = 1'h0;
    440: T381 = 1'h0;
    441: T381 = 1'h0;
    442: T381 = 1'h0;
    443: T381 = 1'h0;
    444: T381 = 1'h0;
    445: T381 = 1'h0;
    446: T381 = 1'h0;
    447: T381 = 1'h0;
    448: T381 = 1'h0;
    449: T381 = 1'h0;
    450: T381 = 1'h0;
    451: T381 = 1'h0;
    452: T381 = 1'h0;
    453: T381 = 1'h0;
    454: T381 = 1'h0;
    455: T381 = 1'h0;
    456: T381 = 1'h0;
    457: T381 = 1'h0;
    458: T381 = 1'h0;
    459: T381 = 1'h0;
    460: T381 = 1'h0;
    461: T381 = 1'h0;
    462: T381 = 1'h0;
    463: T381 = 1'h0;
    464: T381 = 1'h0;
    465: T381 = 1'h0;
    466: T381 = 1'h0;
    467: T381 = 1'h0;
    468: T381 = 1'h0;
    469: T381 = 1'h0;
    470: T381 = 1'h0;
    471: T381 = 1'h0;
    472: T381 = 1'h0;
    473: T381 = 1'h0;
    474: T381 = 1'h0;
    475: T381 = 1'h0;
    476: T381 = 1'h0;
    477: T381 = 1'h0;
    478: T381 = 1'h0;
    479: T381 = 1'h0;
    480: T381 = 1'h0;
    481: T381 = 1'h0;
    482: T381 = 1'h0;
    483: T381 = 1'h0;
    484: T381 = 1'h0;
    485: T381 = 1'h0;
    486: T381 = 1'h0;
    487: T381 = 1'h0;
    488: T381 = 1'h0;
    489: T381 = 1'h0;
    490: T381 = 1'h0;
    491: T381 = 1'h0;
    492: T381 = 1'h0;
    493: T381 = 1'h0;
    494: T381 = 1'h0;
    495: T381 = 1'h0;
    496: T381 = 1'h0;
    497: T381 = 1'h0;
    498: T381 = 1'h0;
    499: T381 = 1'h0;
    500: T381 = 1'h0;
    501: T381 = 1'h0;
    502: T381 = 1'h0;
    503: T381 = 1'h0;
    504: T381 = 1'h0;
    505: T381 = 1'h0;
    506: T381 = 1'h0;
    507: T381 = 1'h0;
    508: T381 = 1'h0;
    509: T381 = 1'h0;
    510: T381 = 1'h0;
    511: T381 = 1'h0;
    512: T381 = 1'h0;
    513: T381 = 1'h0;
    514: T381 = 1'h0;
    515: T381 = 1'h0;
    516: T381 = 1'h0;
    517: T381 = 1'h0;
    518: T381 = 1'h0;
    519: T381 = 1'h0;
    520: T381 = 1'h0;
    521: T381 = 1'h0;
    522: T381 = 1'h0;
    523: T381 = 1'h0;
    524: T381 = 1'h0;
    525: T381 = 1'h0;
    526: T381 = 1'h0;
    527: T381 = 1'h0;
    528: T381 = 1'h0;
    529: T381 = 1'h0;
    530: T381 = 1'h0;
    531: T381 = 1'h0;
    532: T381 = 1'h0;
    533: T381 = 1'h0;
    534: T381 = 1'h0;
    535: T381 = 1'h0;
    536: T381 = 1'h0;
    537: T381 = 1'h0;
    538: T381 = 1'h0;
    539: T381 = 1'h0;
    540: T381 = 1'h0;
    541: T381 = 1'h0;
    542: T381 = 1'h0;
    543: T381 = 1'h0;
    544: T381 = 1'h0;
    545: T381 = 1'h0;
    546: T381 = 1'h0;
    547: T381 = 1'h0;
    548: T381 = 1'h0;
    549: T381 = 1'h0;
    550: T381 = 1'h0;
    551: T381 = 1'h0;
    552: T381 = 1'h0;
    553: T381 = 1'h0;
    554: T381 = 1'h0;
    555: T381 = 1'h0;
    556: T381 = 1'h0;
    557: T381 = 1'h0;
    558: T381 = 1'h0;
    559: T381 = 1'h0;
    560: T381 = 1'h0;
    561: T381 = 1'h0;
    562: T381 = 1'h0;
    563: T381 = 1'h0;
    564: T381 = 1'h0;
    565: T381 = 1'h0;
    566: T381 = 1'h0;
    567: T381 = 1'h0;
    568: T381 = 1'h0;
    569: T381 = 1'h0;
    570: T381 = 1'h0;
    571: T381 = 1'h0;
    572: T381 = 1'h0;
    573: T381 = 1'h0;
    574: T381 = 1'h0;
    575: T381 = 1'h0;
    576: T381 = 1'h0;
    577: T381 = 1'h0;
    578: T381 = 1'h0;
    579: T381 = 1'h0;
    580: T381 = 1'h0;
    581: T381 = 1'h0;
    582: T381 = 1'h0;
    583: T381 = 1'h0;
    584: T381 = 1'h0;
    585: T381 = 1'h0;
    586: T381 = 1'h0;
    587: T381 = 1'h0;
    588: T381 = 1'h0;
    589: T381 = 1'h0;
    590: T381 = 1'h0;
    591: T381 = 1'h0;
    592: T381 = 1'h0;
    593: T381 = 1'h0;
    594: T381 = 1'h0;
    595: T381 = 1'h0;
    596: T381 = 1'h0;
    597: T381 = 1'h0;
    598: T381 = 1'h0;
    599: T381 = 1'h0;
    600: T381 = 1'h0;
    601: T381 = 1'h0;
    602: T381 = 1'h0;
    603: T381 = 1'h0;
    604: T381 = 1'h0;
    605: T381 = 1'h0;
    606: T381 = 1'h0;
    607: T381 = 1'h0;
    608: T381 = 1'h0;
    609: T381 = 1'h0;
    610: T381 = 1'h0;
    611: T381 = 1'h0;
    612: T381 = 1'h0;
    613: T381 = 1'h0;
    614: T381 = 1'h0;
    615: T381 = 1'h0;
    616: T381 = 1'h0;
    617: T381 = 1'h0;
    618: T381 = 1'h0;
    619: T381 = 1'h0;
    620: T381 = 1'h0;
    621: T381 = 1'h0;
    622: T381 = 1'h0;
    623: T381 = 1'h0;
    624: T381 = 1'h0;
    625: T381 = 1'h0;
    626: T381 = 1'h0;
    627: T381 = 1'h0;
    628: T381 = 1'h0;
    629: T381 = 1'h0;
    630: T381 = 1'h0;
    631: T381 = 1'h0;
    632: T381 = 1'h0;
    633: T381 = 1'h0;
    634: T381 = 1'h0;
    635: T381 = 1'h0;
    636: T381 = 1'h0;
    637: T381 = 1'h0;
    638: T381 = 1'h0;
    639: T381 = 1'h0;
    640: T381 = 1'h0;
    641: T381 = 1'h0;
    642: T381 = 1'h0;
    643: T381 = 1'h0;
    644: T381 = 1'h0;
    645: T381 = 1'h0;
    646: T381 = 1'h0;
    647: T381 = 1'h0;
    648: T381 = 1'h0;
    649: T381 = 1'h0;
    650: T381 = 1'h0;
    651: T381 = 1'h0;
    652: T381 = 1'h0;
    653: T381 = 1'h0;
    654: T381 = 1'h0;
    655: T381 = 1'h0;
    656: T381 = 1'h0;
    657: T381 = 1'h0;
    658: T381 = 1'h0;
    659: T381 = 1'h0;
    660: T381 = 1'h0;
    661: T381 = 1'h0;
    662: T381 = 1'h0;
    663: T381 = 1'h0;
    664: T381 = 1'h0;
    665: T381 = 1'h0;
    666: T381 = 1'h0;
    667: T381 = 1'h0;
    668: T381 = 1'h0;
    669: T381 = 1'h0;
    670: T381 = 1'h0;
    671: T381 = 1'h0;
    672: T381 = 1'h0;
    673: T381 = 1'h0;
    674: T381 = 1'h0;
    675: T381 = 1'h0;
    676: T381 = 1'h0;
    677: T381 = 1'h0;
    678: T381 = 1'h0;
    679: T381 = 1'h0;
    680: T381 = 1'h0;
    681: T381 = 1'h0;
    682: T381 = 1'h0;
    683: T381 = 1'h0;
    684: T381 = 1'h0;
    685: T381 = 1'h0;
    686: T381 = 1'h0;
    687: T381 = 1'h0;
    688: T381 = 1'h0;
    689: T381 = 1'h0;
    690: T381 = 1'h0;
    691: T381 = 1'h0;
    692: T381 = 1'h0;
    693: T381 = 1'h0;
    694: T381 = 1'h0;
    695: T381 = 1'h0;
    696: T381 = 1'h0;
    697: T381 = 1'h0;
    698: T381 = 1'h0;
    699: T381 = 1'h0;
    700: T381 = 1'h0;
    701: T381 = 1'h0;
    702: T381 = 1'h0;
    703: T381 = 1'h0;
    704: T381 = 1'h0;
    705: T381 = 1'h0;
    706: T381 = 1'h0;
    707: T381 = 1'h0;
    708: T381 = 1'h0;
    709: T381 = 1'h0;
    710: T381 = 1'h0;
    711: T381 = 1'h0;
    712: T381 = 1'h0;
    713: T381 = 1'h0;
    714: T381 = 1'h0;
    715: T381 = 1'h0;
    716: T381 = 1'h0;
    717: T381 = 1'h0;
    718: T381 = 1'h0;
    719: T381 = 1'h0;
    720: T381 = 1'h0;
    721: T381 = 1'h0;
    722: T381 = 1'h0;
    723: T381 = 1'h0;
    724: T381 = 1'h0;
    725: T381 = 1'h0;
    726: T381 = 1'h0;
    727: T381 = 1'h0;
    728: T381 = 1'h0;
    729: T381 = 1'h0;
    730: T381 = 1'h0;
    731: T381 = 1'h0;
    732: T381 = 1'h0;
    733: T381 = 1'h0;
    734: T381 = 1'h0;
    735: T381 = 1'h0;
    736: T381 = 1'h0;
    737: T381 = 1'h0;
    738: T381 = 1'h0;
    739: T381 = 1'h0;
    740: T381 = 1'h0;
    741: T381 = 1'h0;
    742: T381 = 1'h0;
    743: T381 = 1'h0;
    744: T381 = 1'h0;
    745: T381 = 1'h0;
    746: T381 = 1'h0;
    747: T381 = 1'h0;
    748: T381 = 1'h0;
    749: T381 = 1'h0;
    750: T381 = 1'h0;
    751: T381 = 1'h0;
    752: T381 = 1'h0;
    753: T381 = 1'h0;
    754: T381 = 1'h0;
    755: T381 = 1'h0;
    756: T381 = 1'h0;
    757: T381 = 1'h0;
    758: T381 = 1'h0;
    759: T381 = 1'h0;
    760: T381 = 1'h0;
    761: T381 = 1'h0;
    762: T381 = 1'h0;
    763: T381 = 1'h0;
    764: T381 = 1'h0;
    765: T381 = 1'h0;
    766: T381 = 1'h0;
    767: T381 = 1'h0;
    768: T381 = 1'h0;
    769: T381 = 1'h0;
    770: T381 = 1'h0;
    771: T381 = 1'h0;
    772: T381 = 1'h0;
    773: T381 = 1'h0;
    774: T381 = 1'h0;
    775: T381 = 1'h0;
    776: T381 = 1'h0;
    777: T381 = 1'h0;
    778: T381 = 1'h0;
    779: T381 = 1'h0;
    780: T381 = 1'h0;
    781: T381 = 1'h0;
    782: T381 = 1'h0;
    783: T381 = 1'h0;
    784: T381 = 1'h0;
    785: T381 = 1'h0;
    786: T381 = 1'h0;
    787: T381 = 1'h0;
    788: T381 = 1'h0;
    789: T381 = 1'h0;
    790: T381 = 1'h0;
    791: T381 = 1'h0;
    792: T381 = 1'h0;
    793: T381 = 1'h0;
    794: T381 = 1'h0;
    795: T381 = 1'h0;
    796: T381 = 1'h0;
    797: T381 = 1'h0;
    798: T381 = 1'h0;
    799: T381 = 1'h0;
    800: T381 = 1'h0;
    801: T381 = 1'h0;
    802: T381 = 1'h0;
    803: T381 = 1'h0;
    804: T381 = 1'h0;
    805: T381 = 1'h0;
    806: T381 = 1'h0;
    807: T381 = 1'h0;
    808: T381 = 1'h0;
    809: T381 = 1'h0;
    810: T381 = 1'h0;
    811: T381 = 1'h0;
    812: T381 = 1'h0;
    813: T381 = 1'h0;
    814: T381 = 1'h0;
    815: T381 = 1'h0;
    816: T381 = 1'h0;
    817: T381 = 1'h0;
    818: T381 = 1'h0;
    819: T381 = 1'h0;
    820: T381 = 1'h0;
    821: T381 = 1'h0;
    822: T381 = 1'h0;
    823: T381 = 1'h0;
    824: T381 = 1'h0;
    825: T381 = 1'h0;
    826: T381 = 1'h0;
    827: T381 = 1'h0;
    828: T381 = 1'h0;
    829: T381 = 1'h0;
    830: T381 = 1'h0;
    831: T381 = 1'h0;
    832: T381 = 1'h0;
    833: T381 = 1'h0;
    834: T381 = 1'h0;
    835: T381 = 1'h0;
    836: T381 = 1'h0;
    837: T381 = 1'h0;
    838: T381 = 1'h0;
    839: T381 = 1'h0;
    840: T381 = 1'h0;
    841: T381 = 1'h0;
    842: T381 = 1'h0;
    843: T381 = 1'h0;
    844: T381 = 1'h0;
    845: T381 = 1'h0;
    846: T381 = 1'h0;
    847: T381 = 1'h0;
    848: T381 = 1'h0;
    849: T381 = 1'h0;
    850: T381 = 1'h0;
    851: T381 = 1'h0;
    852: T381 = 1'h0;
    853: T381 = 1'h0;
    854: T381 = 1'h0;
    855: T381 = 1'h0;
    856: T381 = 1'h0;
    857: T381 = 1'h0;
    858: T381 = 1'h0;
    859: T381 = 1'h0;
    860: T381 = 1'h0;
    861: T381 = 1'h0;
    862: T381 = 1'h0;
    863: T381 = 1'h0;
    864: T381 = 1'h0;
    865: T381 = 1'h0;
    866: T381 = 1'h0;
    867: T381 = 1'h0;
    868: T381 = 1'h0;
    869: T381 = 1'h0;
    870: T381 = 1'h0;
    871: T381 = 1'h0;
    872: T381 = 1'h0;
    873: T381 = 1'h0;
    874: T381 = 1'h0;
    875: T381 = 1'h0;
    876: T381 = 1'h0;
    877: T381 = 1'h0;
    878: T381 = 1'h0;
    879: T381 = 1'h0;
    880: T381 = 1'h0;
    881: T381 = 1'h0;
    882: T381 = 1'h0;
    883: T381 = 1'h0;
    884: T381 = 1'h0;
    885: T381 = 1'h0;
    886: T381 = 1'h0;
    887: T381 = 1'h0;
    888: T381 = 1'h0;
    889: T381 = 1'h0;
    890: T381 = 1'h0;
    891: T381 = 1'h0;
    892: T381 = 1'h0;
    893: T381 = 1'h0;
    894: T381 = 1'h0;
    895: T381 = 1'h0;
    896: T381 = 1'h0;
    897: T381 = 1'h0;
    898: T381 = 1'h0;
    899: T381 = 1'h0;
    900: T381 = 1'h0;
    901: T381 = 1'h0;
    902: T381 = 1'h0;
    903: T381 = 1'h0;
    904: T381 = 1'h0;
    905: T381 = 1'h0;
    906: T381 = 1'h0;
    907: T381 = 1'h0;
    908: T381 = 1'h0;
    909: T381 = 1'h0;
    910: T381 = 1'h0;
    911: T381 = 1'h0;
    912: T381 = 1'h0;
    913: T381 = 1'h0;
    914: T381 = 1'h0;
    915: T381 = 1'h0;
    916: T381 = 1'h0;
    917: T381 = 1'h0;
    918: T381 = 1'h0;
    919: T381 = 1'h0;
    920: T381 = 1'h0;
    921: T381 = 1'h0;
    922: T381 = 1'h0;
    923: T381 = 1'h0;
    924: T381 = 1'h0;
    925: T381 = 1'h0;
    926: T381 = 1'h0;
    927: T381 = 1'h0;
    928: T381 = 1'h0;
    929: T381 = 1'h0;
    930: T381 = 1'h0;
    931: T381 = 1'h0;
    932: T381 = 1'h0;
    933: T381 = 1'h0;
    934: T381 = 1'h0;
    935: T381 = 1'h0;
    936: T381 = 1'h0;
    937: T381 = 1'h0;
    938: T381 = 1'h0;
    939: T381 = 1'h0;
    940: T381 = 1'h0;
    941: T381 = 1'h0;
    942: T381 = 1'h0;
    943: T381 = 1'h0;
    944: T381 = 1'h0;
    945: T381 = 1'h0;
    946: T381 = 1'h0;
    947: T381 = 1'h0;
    948: T381 = 1'h0;
    949: T381 = 1'h0;
    950: T381 = 1'h0;
    951: T381 = 1'h0;
    952: T381 = 1'h0;
    953: T381 = 1'h0;
    954: T381 = 1'h0;
    955: T381 = 1'h0;
    956: T381 = 1'h0;
    957: T381 = 1'h0;
    958: T381 = 1'h0;
    959: T381 = 1'h0;
    960: T381 = 1'h0;
    961: T381 = 1'h0;
    962: T381 = 1'h0;
    963: T381 = 1'h0;
    964: T381 = 1'h0;
    965: T381 = 1'h0;
    966: T381 = 1'h0;
    967: T381 = 1'h0;
    968: T381 = 1'h0;
    969: T381 = 1'h0;
    970: T381 = 1'h0;
    971: T381 = 1'h0;
    972: T381 = 1'h0;
    973: T381 = 1'h0;
    974: T381 = 1'h0;
    975: T381 = 1'h0;
    976: T381 = 1'h0;
    977: T381 = 1'h0;
    978: T381 = 1'h0;
    979: T381 = 1'h0;
    980: T381 = 1'h0;
    981: T381 = 1'h0;
    982: T381 = 1'h0;
    983: T381 = 1'h0;
    984: T381 = 1'h0;
    985: T381 = 1'h0;
    986: T381 = 1'h0;
    987: T381 = 1'h0;
    988: T381 = 1'h0;
    989: T381 = 1'h0;
    990: T381 = 1'h0;
    991: T381 = 1'h0;
    992: T381 = 1'h0;
    993: T381 = 1'h0;
    994: T381 = 1'h0;
    995: T381 = 1'h0;
    996: T381 = 1'h0;
    997: T381 = 1'h0;
    998: T381 = 1'h0;
    999: T381 = 1'h0;
    1000: T381 = 1'h0;
    1001: T381 = 1'h0;
    1002: T381 = 1'h0;
    1003: T381 = 1'h0;
    1004: T381 = 1'h0;
    1005: T381 = 1'h0;
    1006: T381 = 1'h0;
    1007: T381 = 1'h0;
    1008: T381 = 1'h0;
    1009: T381 = 1'h0;
    1010: T381 = 1'h0;
    1011: T381 = 1'h0;
    1012: T381 = 1'h0;
    1013: T381 = 1'h0;
    1014: T381 = 1'h0;
    1015: T381 = 1'h0;
    1016: T381 = 1'h0;
    1017: T381 = 1'h0;
    1018: T381 = 1'h0;
    1019: T381 = 1'h0;
    1020: T381 = 1'h0;
    1021: T381 = 1'h0;
    1022: T381 = 1'h0;
    1023: T381 = 1'h0;
    1024: T381 = 1'h0;
    1025: T381 = 1'h0;
    1026: T381 = 1'h0;
    1027: T381 = 1'h0;
    1028: T381 = 1'h0;
    1029: T381 = 1'h0;
    1030: T381 = 1'h0;
    1031: T381 = 1'h0;
    1032: T381 = 1'h0;
    1033: T381 = 1'h0;
    1034: T381 = 1'h0;
    1035: T381 = 1'h0;
    1036: T381 = 1'h0;
    1037: T381 = 1'h0;
    1038: T381 = 1'h0;
    1039: T381 = 1'h0;
    1040: T381 = 1'h0;
    1041: T381 = 1'h0;
    1042: T381 = 1'h0;
    1043: T381 = 1'h0;
    1044: T381 = 1'h0;
    1045: T381 = 1'h0;
    1046: T381 = 1'h0;
    1047: T381 = 1'h0;
    1048: T381 = 1'h0;
    1049: T381 = 1'h0;
    1050: T381 = 1'h0;
    1051: T381 = 1'h0;
    1052: T381 = 1'h0;
    1053: T381 = 1'h0;
    1054: T381 = 1'h0;
    1055: T381 = 1'h0;
    1056: T381 = 1'h0;
    1057: T381 = 1'h0;
    1058: T381 = 1'h0;
    1059: T381 = 1'h0;
    1060: T381 = 1'h0;
    1061: T381 = 1'h0;
    1062: T381 = 1'h0;
    1063: T381 = 1'h0;
    1064: T381 = 1'h0;
    1065: T381 = 1'h0;
    1066: T381 = 1'h0;
    1067: T381 = 1'h0;
    1068: T381 = 1'h0;
    1069: T381 = 1'h0;
    1070: T381 = 1'h0;
    1071: T381 = 1'h0;
    1072: T381 = 1'h0;
    1073: T381 = 1'h0;
    1074: T381 = 1'h0;
    1075: T381 = 1'h0;
    1076: T381 = 1'h0;
    1077: T381 = 1'h0;
    1078: T381 = 1'h0;
    1079: T381 = 1'h0;
    1080: T381 = 1'h0;
    1081: T381 = 1'h0;
    1082: T381 = 1'h0;
    1083: T381 = 1'h0;
    1084: T381 = 1'h0;
    1085: T381 = 1'h0;
    1086: T381 = 1'h0;
    1087: T381 = 1'h0;
    1088: T381 = 1'h0;
    1089: T381 = 1'h0;
    1090: T381 = 1'h0;
    1091: T381 = 1'h0;
    1092: T381 = 1'h0;
    1093: T381 = 1'h0;
    1094: T381 = 1'h0;
    1095: T381 = 1'h0;
    1096: T381 = 1'h0;
    1097: T381 = 1'h0;
    1098: T381 = 1'h0;
    1099: T381 = 1'h0;
    1100: T381 = 1'h0;
    1101: T381 = 1'h0;
    1102: T381 = 1'h0;
    1103: T381 = 1'h0;
    1104: T381 = 1'h0;
    1105: T381 = 1'h0;
    1106: T381 = 1'h0;
    1107: T381 = 1'h0;
    1108: T381 = 1'h0;
    1109: T381 = 1'h0;
    1110: T381 = 1'h0;
    1111: T381 = 1'h0;
    1112: T381 = 1'h0;
    1113: T381 = 1'h0;
    1114: T381 = 1'h0;
    1115: T381 = 1'h0;
    1116: T381 = 1'h0;
    1117: T381 = 1'h0;
    1118: T381 = 1'h0;
    1119: T381 = 1'h0;
    1120: T381 = 1'h0;
    1121: T381 = 1'h0;
    1122: T381 = 1'h0;
    1123: T381 = 1'h0;
    1124: T381 = 1'h0;
    1125: T381 = 1'h0;
    1126: T381 = 1'h0;
    1127: T381 = 1'h0;
    1128: T381 = 1'h0;
    1129: T381 = 1'h0;
    1130: T381 = 1'h0;
    1131: T381 = 1'h0;
    1132: T381 = 1'h0;
    1133: T381 = 1'h0;
    1134: T381 = 1'h0;
    1135: T381 = 1'h0;
    1136: T381 = 1'h0;
    1137: T381 = 1'h0;
    1138: T381 = 1'h0;
    1139: T381 = 1'h0;
    1140: T381 = 1'h0;
    1141: T381 = 1'h0;
    1142: T381 = 1'h0;
    1143: T381 = 1'h0;
    1144: T381 = 1'h0;
    1145: T381 = 1'h0;
    1146: T381 = 1'h0;
    1147: T381 = 1'h0;
    1148: T381 = 1'h0;
    1149: T381 = 1'h0;
    1150: T381 = 1'h0;
    1151: T381 = 1'h0;
    1152: T381 = 1'h0;
    1153: T381 = 1'h0;
    1154: T381 = 1'h0;
    1155: T381 = 1'h0;
    1156: T381 = 1'h0;
    1157: T381 = 1'h0;
    1158: T381 = 1'h0;
    1159: T381 = 1'h0;
    1160: T381 = 1'h0;
    1161: T381 = 1'h0;
    1162: T381 = 1'h0;
    1163: T381 = 1'h0;
    1164: T381 = 1'h0;
    1165: T381 = 1'h0;
    1166: T381 = 1'h0;
    1167: T381 = 1'h0;
    1168: T381 = 1'h0;
    1169: T381 = 1'h0;
    1170: T381 = 1'h0;
    1171: T381 = 1'h0;
    1172: T381 = 1'h0;
    1173: T381 = 1'h0;
    1174: T381 = 1'h0;
    1175: T381 = 1'h0;
    1176: T381 = 1'h0;
    1177: T381 = 1'h0;
    1178: T381 = 1'h0;
    1179: T381 = 1'h0;
    1180: T381 = 1'h0;
    1181: T381 = 1'h0;
    1182: T381 = 1'h0;
    1183: T381 = 1'h0;
    1184: T381 = 1'h0;
    1185: T381 = 1'h0;
    1186: T381 = 1'h0;
    1187: T381 = 1'h0;
    1188: T381 = 1'h0;
    1189: T381 = 1'h0;
    1190: T381 = 1'h0;
    1191: T381 = 1'h0;
    1192: T381 = 1'h0;
    1193: T381 = 1'h0;
    1194: T381 = 1'h0;
    1195: T381 = 1'h0;
    1196: T381 = 1'h0;
    1197: T381 = 1'h0;
    1198: T381 = 1'h0;
    1199: T381 = 1'h0;
    1200: T381 = 1'h0;
    1201: T381 = 1'h0;
    1202: T381 = 1'h0;
    1203: T381 = 1'h0;
    1204: T381 = 1'h0;
    1205: T381 = 1'h0;
    1206: T381 = 1'h0;
    1207: T381 = 1'h0;
    1208: T381 = 1'h0;
    1209: T381 = 1'h0;
    1210: T381 = 1'h0;
    1211: T381 = 1'h0;
    1212: T381 = 1'h0;
    1213: T381 = 1'h0;
    1214: T381 = 1'h0;
    1215: T381 = 1'h0;
    1216: T381 = 1'h0;
    1217: T381 = 1'h0;
    1218: T381 = 1'h0;
    1219: T381 = 1'h0;
    1220: T381 = 1'h0;
    1221: T381 = 1'h0;
    1222: T381 = 1'h0;
    1223: T381 = 1'h0;
    1224: T381 = 1'h0;
    1225: T381 = 1'h0;
    1226: T381 = 1'h0;
    1227: T381 = 1'h0;
    1228: T381 = 1'h0;
    1229: T381 = 1'h0;
    1230: T381 = 1'h0;
    1231: T381 = 1'h0;
    1232: T381 = 1'h0;
    1233: T381 = 1'h0;
    1234: T381 = 1'h0;
    1235: T381 = 1'h0;
    1236: T381 = 1'h0;
    1237: T381 = 1'h0;
    1238: T381 = 1'h0;
    1239: T381 = 1'h0;
    1240: T381 = 1'h0;
    1241: T381 = 1'h0;
    1242: T381 = 1'h0;
    1243: T381 = 1'h0;
    1244: T381 = 1'h0;
    1245: T381 = 1'h0;
    1246: T381 = 1'h0;
    1247: T381 = 1'h0;
    1248: T381 = 1'h0;
    1249: T381 = 1'h0;
    1250: T381 = 1'h0;
    1251: T381 = 1'h0;
    1252: T381 = 1'h0;
    1253: T381 = 1'h0;
    1254: T381 = 1'h0;
    1255: T381 = 1'h0;
    1256: T381 = 1'h0;
    1257: T381 = 1'h0;
    1258: T381 = 1'h0;
    1259: T381 = 1'h0;
    1260: T381 = 1'h0;
    1261: T381 = 1'h0;
    1262: T381 = 1'h0;
    1263: T381 = 1'h0;
    1264: T381 = 1'h0;
    1265: T381 = 1'h0;
    1266: T381 = 1'h0;
    1267: T381 = 1'h0;
    1268: T381 = 1'h0;
    1269: T381 = 1'h0;
    1270: T381 = 1'h0;
    1271: T381 = 1'h0;
    1272: T381 = 1'h0;
    1273: T381 = 1'h0;
    1274: T381 = 1'h0;
    1275: T381 = 1'h0;
    1276: T381 = 1'h0;
    1277: T381 = 1'h0;
    1278: T381 = 1'h0;
    1279: T381 = 1'h0;
    1280: T381 = 1'h1;
    1281: T381 = 1'h1;
    1282: T381 = 1'h1;
    1283: T381 = 1'h1;
    1284: T381 = 1'h1;
    1285: T381 = 1'h1;
    1286: T381 = 1'h1;
    1287: T381 = 1'h1;
    1288: T381 = 1'h1;
    1289: T381 = 1'h1;
    1290: T381 = 1'h1;
    1291: T381 = 1'h1;
    1292: T381 = 1'h1;
    1293: T381 = 1'h1;
    1294: T381 = 1'h1;
    1295: T381 = 1'h1;
    1296: T381 = 1'h0;
    1297: T381 = 1'h0;
    1298: T381 = 1'h0;
    1299: T381 = 1'h0;
    1300: T381 = 1'h0;
    1301: T381 = 1'h0;
    1302: T381 = 1'h0;
    1303: T381 = 1'h0;
    1304: T381 = 1'h0;
    1305: T381 = 1'h0;
    1306: T381 = 1'h0;
    1307: T381 = 1'h0;
    1308: T381 = 1'h0;
    1309: T381 = 1'h1;
    1310: T381 = 1'h1;
    1311: T381 = 1'h1;
    1312: T381 = 1'h0;
    1313: T381 = 1'h0;
    1314: T381 = 1'h0;
    1315: T381 = 1'h0;
    1316: T381 = 1'h0;
    1317: T381 = 1'h0;
    1318: T381 = 1'h0;
    1319: T381 = 1'h0;
    1320: T381 = 1'h0;
    1321: T381 = 1'h0;
    1322: T381 = 1'h0;
    1323: T381 = 1'h0;
    1324: T381 = 1'h0;
    1325: T381 = 1'h0;
    1326: T381 = 1'h0;
    1327: T381 = 1'h0;
    1328: T381 = 1'h0;
    1329: T381 = 1'h0;
    1330: T381 = 1'h0;
    1331: T381 = 1'h0;
    1332: T381 = 1'h0;
    1333: T381 = 1'h0;
    1334: T381 = 1'h0;
    1335: T381 = 1'h0;
    1336: T381 = 1'h0;
    1337: T381 = 1'h0;
    1338: T381 = 1'h0;
    1339: T381 = 1'h0;
    1340: T381 = 1'h0;
    1341: T381 = 1'h0;
    1342: T381 = 1'h0;
    1343: T381 = 1'h0;
    1344: T381 = 1'h0;
    1345: T381 = 1'h0;
    1346: T381 = 1'h0;
    1347: T381 = 1'h0;
    1348: T381 = 1'h0;
    1349: T381 = 1'h0;
    1350: T381 = 1'h0;
    1351: T381 = 1'h0;
    1352: T381 = 1'h0;
    1353: T381 = 1'h0;
    1354: T381 = 1'h0;
    1355: T381 = 1'h0;
    1356: T381 = 1'h0;
    1357: T381 = 1'h0;
    1358: T381 = 1'h0;
    1359: T381 = 1'h0;
    1360: T381 = 1'h0;
    1361: T381 = 1'h0;
    1362: T381 = 1'h0;
    1363: T381 = 1'h0;
    1364: T381 = 1'h0;
    1365: T381 = 1'h0;
    1366: T381 = 1'h0;
    1367: T381 = 1'h0;
    1368: T381 = 1'h0;
    1369: T381 = 1'h0;
    1370: T381 = 1'h0;
    1371: T381 = 1'h0;
    1372: T381 = 1'h0;
    1373: T381 = 1'h0;
    1374: T381 = 1'h0;
    1375: T381 = 1'h0;
    1376: T381 = 1'h0;
    1377: T381 = 1'h0;
    1378: T381 = 1'h0;
    1379: T381 = 1'h0;
    1380: T381 = 1'h0;
    1381: T381 = 1'h0;
    1382: T381 = 1'h0;
    1383: T381 = 1'h0;
    1384: T381 = 1'h0;
    1385: T381 = 1'h0;
    1386: T381 = 1'h0;
    1387: T381 = 1'h0;
    1388: T381 = 1'h0;
    1389: T381 = 1'h0;
    1390: T381 = 1'h0;
    1391: T381 = 1'h0;
    1392: T381 = 1'h0;
    1393: T381 = 1'h0;
    1394: T381 = 1'h0;
    1395: T381 = 1'h0;
    1396: T381 = 1'h0;
    1397: T381 = 1'h0;
    1398: T381 = 1'h0;
    1399: T381 = 1'h0;
    1400: T381 = 1'h0;
    1401: T381 = 1'h0;
    1402: T381 = 1'h0;
    1403: T381 = 1'h0;
    1404: T381 = 1'h0;
    1405: T381 = 1'h0;
    1406: T381 = 1'h0;
    1407: T381 = 1'h0;
    1408: T381 = 1'h0;
    1409: T381 = 1'h0;
    1410: T381 = 1'h0;
    1411: T381 = 1'h0;
    1412: T381 = 1'h0;
    1413: T381 = 1'h0;
    1414: T381 = 1'h0;
    1415: T381 = 1'h0;
    1416: T381 = 1'h0;
    1417: T381 = 1'h0;
    1418: T381 = 1'h0;
    1419: T381 = 1'h0;
    1420: T381 = 1'h0;
    1421: T381 = 1'h0;
    1422: T381 = 1'h0;
    1423: T381 = 1'h0;
    1424: T381 = 1'h0;
    1425: T381 = 1'h0;
    1426: T381 = 1'h0;
    1427: T381 = 1'h0;
    1428: T381 = 1'h0;
    1429: T381 = 1'h0;
    1430: T381 = 1'h0;
    1431: T381 = 1'h0;
    1432: T381 = 1'h0;
    1433: T381 = 1'h0;
    1434: T381 = 1'h0;
    1435: T381 = 1'h0;
    1436: T381 = 1'h0;
    1437: T381 = 1'h0;
    1438: T381 = 1'h0;
    1439: T381 = 1'h0;
    1440: T381 = 1'h0;
    1441: T381 = 1'h0;
    1442: T381 = 1'h0;
    1443: T381 = 1'h0;
    1444: T381 = 1'h0;
    1445: T381 = 1'h0;
    1446: T381 = 1'h0;
    1447: T381 = 1'h0;
    1448: T381 = 1'h0;
    1449: T381 = 1'h0;
    1450: T381 = 1'h0;
    1451: T381 = 1'h0;
    1452: T381 = 1'h0;
    1453: T381 = 1'h0;
    1454: T381 = 1'h0;
    1455: T381 = 1'h0;
    1456: T381 = 1'h0;
    1457: T381 = 1'h0;
    1458: T381 = 1'h0;
    1459: T381 = 1'h0;
    1460: T381 = 1'h0;
    1461: T381 = 1'h0;
    1462: T381 = 1'h0;
    1463: T381 = 1'h0;
    1464: T381 = 1'h0;
    1465: T381 = 1'h0;
    1466: T381 = 1'h0;
    1467: T381 = 1'h0;
    1468: T381 = 1'h0;
    1469: T381 = 1'h0;
    1470: T381 = 1'h0;
    1471: T381 = 1'h0;
    1472: T381 = 1'h0;
    1473: T381 = 1'h0;
    1474: T381 = 1'h0;
    1475: T381 = 1'h0;
    1476: T381 = 1'h0;
    1477: T381 = 1'h0;
    1478: T381 = 1'h0;
    1479: T381 = 1'h0;
    1480: T381 = 1'h0;
    1481: T381 = 1'h0;
    1482: T381 = 1'h0;
    1483: T381 = 1'h0;
    1484: T381 = 1'h0;
    1485: T381 = 1'h0;
    1486: T381 = 1'h0;
    1487: T381 = 1'h0;
    1488: T381 = 1'h0;
    1489: T381 = 1'h0;
    1490: T381 = 1'h0;
    1491: T381 = 1'h0;
    1492: T381 = 1'h0;
    1493: T381 = 1'h0;
    1494: T381 = 1'h0;
    1495: T381 = 1'h0;
    1496: T381 = 1'h0;
    1497: T381 = 1'h0;
    1498: T381 = 1'h0;
    1499: T381 = 1'h0;
    1500: T381 = 1'h0;
    1501: T381 = 1'h0;
    1502: T381 = 1'h0;
    1503: T381 = 1'h0;
    1504: T381 = 1'h0;
    1505: T381 = 1'h0;
    1506: T381 = 1'h0;
    1507: T381 = 1'h0;
    1508: T381 = 1'h0;
    1509: T381 = 1'h0;
    1510: T381 = 1'h0;
    1511: T381 = 1'h0;
    1512: T381 = 1'h0;
    1513: T381 = 1'h0;
    1514: T381 = 1'h0;
    1515: T381 = 1'h0;
    1516: T381 = 1'h0;
    1517: T381 = 1'h0;
    1518: T381 = 1'h0;
    1519: T381 = 1'h0;
    1520: T381 = 1'h0;
    1521: T381 = 1'h0;
    1522: T381 = 1'h0;
    1523: T381 = 1'h0;
    1524: T381 = 1'h0;
    1525: T381 = 1'h0;
    1526: T381 = 1'h0;
    1527: T381 = 1'h0;
    1528: T381 = 1'h0;
    1529: T381 = 1'h0;
    1530: T381 = 1'h0;
    1531: T381 = 1'h0;
    1532: T381 = 1'h0;
    1533: T381 = 1'h0;
    1534: T381 = 1'h0;
    1535: T381 = 1'h0;
    1536: T381 = 1'h0;
    1537: T381 = 1'h0;
    1538: T381 = 1'h0;
    1539: T381 = 1'h0;
    1540: T381 = 1'h0;
    1541: T381 = 1'h0;
    1542: T381 = 1'h0;
    1543: T381 = 1'h0;
    1544: T381 = 1'h0;
    1545: T381 = 1'h0;
    1546: T381 = 1'h0;
    1547: T381 = 1'h0;
    1548: T381 = 1'h0;
    1549: T381 = 1'h0;
    1550: T381 = 1'h0;
    1551: T381 = 1'h0;
    1552: T381 = 1'h0;
    1553: T381 = 1'h0;
    1554: T381 = 1'h0;
    1555: T381 = 1'h0;
    1556: T381 = 1'h0;
    1557: T381 = 1'h0;
    1558: T381 = 1'h0;
    1559: T381 = 1'h0;
    1560: T381 = 1'h0;
    1561: T381 = 1'h0;
    1562: T381 = 1'h0;
    1563: T381 = 1'h0;
    1564: T381 = 1'h0;
    1565: T381 = 1'h0;
    1566: T381 = 1'h0;
    1567: T381 = 1'h0;
    1568: T381 = 1'h0;
    1569: T381 = 1'h0;
    1570: T381 = 1'h0;
    1571: T381 = 1'h0;
    1572: T381 = 1'h0;
    1573: T381 = 1'h0;
    1574: T381 = 1'h0;
    1575: T381 = 1'h0;
    1576: T381 = 1'h0;
    1577: T381 = 1'h0;
    1578: T381 = 1'h0;
    1579: T381 = 1'h0;
    1580: T381 = 1'h0;
    1581: T381 = 1'h0;
    1582: T381 = 1'h0;
    1583: T381 = 1'h0;
    1584: T381 = 1'h0;
    1585: T381 = 1'h0;
    1586: T381 = 1'h0;
    1587: T381 = 1'h0;
    1588: T381 = 1'h0;
    1589: T381 = 1'h0;
    1590: T381 = 1'h0;
    1591: T381 = 1'h0;
    1592: T381 = 1'h0;
    1593: T381 = 1'h0;
    1594: T381 = 1'h0;
    1595: T381 = 1'h0;
    1596: T381 = 1'h0;
    1597: T381 = 1'h0;
    1598: T381 = 1'h0;
    1599: T381 = 1'h0;
    1600: T381 = 1'h0;
    1601: T381 = 1'h0;
    1602: T381 = 1'h0;
    1603: T381 = 1'h0;
    1604: T381 = 1'h0;
    1605: T381 = 1'h0;
    1606: T381 = 1'h0;
    1607: T381 = 1'h0;
    1608: T381 = 1'h0;
    1609: T381 = 1'h0;
    1610: T381 = 1'h0;
    1611: T381 = 1'h0;
    1612: T381 = 1'h0;
    1613: T381 = 1'h0;
    1614: T381 = 1'h0;
    1615: T381 = 1'h0;
    1616: T381 = 1'h0;
    1617: T381 = 1'h0;
    1618: T381 = 1'h0;
    1619: T381 = 1'h0;
    1620: T381 = 1'h0;
    1621: T381 = 1'h0;
    1622: T381 = 1'h0;
    1623: T381 = 1'h0;
    1624: T381 = 1'h0;
    1625: T381 = 1'h0;
    1626: T381 = 1'h0;
    1627: T381 = 1'h0;
    1628: T381 = 1'h0;
    1629: T381 = 1'h0;
    1630: T381 = 1'h0;
    1631: T381 = 1'h0;
    1632: T381 = 1'h0;
    1633: T381 = 1'h0;
    1634: T381 = 1'h0;
    1635: T381 = 1'h0;
    1636: T381 = 1'h0;
    1637: T381 = 1'h0;
    1638: T381 = 1'h0;
    1639: T381 = 1'h0;
    1640: T381 = 1'h0;
    1641: T381 = 1'h0;
    1642: T381 = 1'h0;
    1643: T381 = 1'h0;
    1644: T381 = 1'h0;
    1645: T381 = 1'h0;
    1646: T381 = 1'h0;
    1647: T381 = 1'h0;
    1648: T381 = 1'h0;
    1649: T381 = 1'h0;
    1650: T381 = 1'h0;
    1651: T381 = 1'h0;
    1652: T381 = 1'h0;
    1653: T381 = 1'h0;
    1654: T381 = 1'h0;
    1655: T381 = 1'h0;
    1656: T381 = 1'h0;
    1657: T381 = 1'h0;
    1658: T381 = 1'h0;
    1659: T381 = 1'h0;
    1660: T381 = 1'h0;
    1661: T381 = 1'h0;
    1662: T381 = 1'h0;
    1663: T381 = 1'h0;
    1664: T381 = 1'h0;
    1665: T381 = 1'h0;
    1666: T381 = 1'h0;
    1667: T381 = 1'h0;
    1668: T381 = 1'h0;
    1669: T381 = 1'h0;
    1670: T381 = 1'h0;
    1671: T381 = 1'h0;
    1672: T381 = 1'h0;
    1673: T381 = 1'h0;
    1674: T381 = 1'h0;
    1675: T381 = 1'h0;
    1676: T381 = 1'h0;
    1677: T381 = 1'h0;
    1678: T381 = 1'h0;
    1679: T381 = 1'h0;
    1680: T381 = 1'h0;
    1681: T381 = 1'h0;
    1682: T381 = 1'h0;
    1683: T381 = 1'h0;
    1684: T381 = 1'h0;
    1685: T381 = 1'h0;
    1686: T381 = 1'h0;
    1687: T381 = 1'h0;
    1688: T381 = 1'h0;
    1689: T381 = 1'h0;
    1690: T381 = 1'h0;
    1691: T381 = 1'h0;
    1692: T381 = 1'h0;
    1693: T381 = 1'h0;
    1694: T381 = 1'h0;
    1695: T381 = 1'h0;
    1696: T381 = 1'h0;
    1697: T381 = 1'h0;
    1698: T381 = 1'h0;
    1699: T381 = 1'h0;
    1700: T381 = 1'h0;
    1701: T381 = 1'h0;
    1702: T381 = 1'h0;
    1703: T381 = 1'h0;
    1704: T381 = 1'h0;
    1705: T381 = 1'h0;
    1706: T381 = 1'h0;
    1707: T381 = 1'h0;
    1708: T381 = 1'h0;
    1709: T381 = 1'h0;
    1710: T381 = 1'h0;
    1711: T381 = 1'h0;
    1712: T381 = 1'h0;
    1713: T381 = 1'h0;
    1714: T381 = 1'h0;
    1715: T381 = 1'h0;
    1716: T381 = 1'h0;
    1717: T381 = 1'h0;
    1718: T381 = 1'h0;
    1719: T381 = 1'h0;
    1720: T381 = 1'h0;
    1721: T381 = 1'h0;
    1722: T381 = 1'h0;
    1723: T381 = 1'h0;
    1724: T381 = 1'h0;
    1725: T381 = 1'h0;
    1726: T381 = 1'h0;
    1727: T381 = 1'h0;
    1728: T381 = 1'h0;
    1729: T381 = 1'h0;
    1730: T381 = 1'h0;
    1731: T381 = 1'h0;
    1732: T381 = 1'h0;
    1733: T381 = 1'h0;
    1734: T381 = 1'h0;
    1735: T381 = 1'h0;
    1736: T381 = 1'h0;
    1737: T381 = 1'h0;
    1738: T381 = 1'h0;
    1739: T381 = 1'h0;
    1740: T381 = 1'h0;
    1741: T381 = 1'h0;
    1742: T381 = 1'h0;
    1743: T381 = 1'h0;
    1744: T381 = 1'h0;
    1745: T381 = 1'h0;
    1746: T381 = 1'h0;
    1747: T381 = 1'h0;
    1748: T381 = 1'h0;
    1749: T381 = 1'h0;
    1750: T381 = 1'h0;
    1751: T381 = 1'h0;
    1752: T381 = 1'h0;
    1753: T381 = 1'h0;
    1754: T381 = 1'h0;
    1755: T381 = 1'h0;
    1756: T381 = 1'h0;
    1757: T381 = 1'h0;
    1758: T381 = 1'h0;
    1759: T381 = 1'h0;
    1760: T381 = 1'h0;
    1761: T381 = 1'h0;
    1762: T381 = 1'h0;
    1763: T381 = 1'h0;
    1764: T381 = 1'h0;
    1765: T381 = 1'h0;
    1766: T381 = 1'h0;
    1767: T381 = 1'h0;
    1768: T381 = 1'h0;
    1769: T381 = 1'h0;
    1770: T381 = 1'h0;
    1771: T381 = 1'h0;
    1772: T381 = 1'h0;
    1773: T381 = 1'h0;
    1774: T381 = 1'h0;
    1775: T381 = 1'h0;
    1776: T381 = 1'h0;
    1777: T381 = 1'h0;
    1778: T381 = 1'h0;
    1779: T381 = 1'h0;
    1780: T381 = 1'h0;
    1781: T381 = 1'h0;
    1782: T381 = 1'h0;
    1783: T381 = 1'h0;
    1784: T381 = 1'h0;
    1785: T381 = 1'h0;
    1786: T381 = 1'h0;
    1787: T381 = 1'h0;
    1788: T381 = 1'h0;
    1789: T381 = 1'h0;
    1790: T381 = 1'h0;
    1791: T381 = 1'h0;
    1792: T381 = 1'h0;
    1793: T381 = 1'h0;
    1794: T381 = 1'h0;
    1795: T381 = 1'h0;
    1796: T381 = 1'h0;
    1797: T381 = 1'h0;
    1798: T381 = 1'h0;
    1799: T381 = 1'h0;
    1800: T381 = 1'h0;
    1801: T381 = 1'h0;
    1802: T381 = 1'h0;
    1803: T381 = 1'h0;
    1804: T381 = 1'h0;
    1805: T381 = 1'h0;
    1806: T381 = 1'h0;
    1807: T381 = 1'h0;
    1808: T381 = 1'h0;
    1809: T381 = 1'h0;
    1810: T381 = 1'h0;
    1811: T381 = 1'h0;
    1812: T381 = 1'h0;
    1813: T381 = 1'h0;
    1814: T381 = 1'h0;
    1815: T381 = 1'h0;
    1816: T381 = 1'h0;
    1817: T381 = 1'h0;
    1818: T381 = 1'h0;
    1819: T381 = 1'h0;
    1820: T381 = 1'h0;
    1821: T381 = 1'h0;
    1822: T381 = 1'h0;
    1823: T381 = 1'h0;
    1824: T381 = 1'h0;
    1825: T381 = 1'h0;
    1826: T381 = 1'h0;
    1827: T381 = 1'h0;
    1828: T381 = 1'h0;
    1829: T381 = 1'h0;
    1830: T381 = 1'h0;
    1831: T381 = 1'h0;
    1832: T381 = 1'h0;
    1833: T381 = 1'h0;
    1834: T381 = 1'h0;
    1835: T381 = 1'h0;
    1836: T381 = 1'h0;
    1837: T381 = 1'h0;
    1838: T381 = 1'h0;
    1839: T381 = 1'h0;
    1840: T381 = 1'h0;
    1841: T381 = 1'h0;
    1842: T381 = 1'h0;
    1843: T381 = 1'h0;
    1844: T381 = 1'h0;
    1845: T381 = 1'h0;
    1846: T381 = 1'h0;
    1847: T381 = 1'h0;
    1848: T381 = 1'h0;
    1849: T381 = 1'h0;
    1850: T381 = 1'h0;
    1851: T381 = 1'h0;
    1852: T381 = 1'h0;
    1853: T381 = 1'h0;
    1854: T381 = 1'h0;
    1855: T381 = 1'h0;
    1856: T381 = 1'h0;
    1857: T381 = 1'h0;
    1858: T381 = 1'h0;
    1859: T381 = 1'h0;
    1860: T381 = 1'h0;
    1861: T381 = 1'h0;
    1862: T381 = 1'h0;
    1863: T381 = 1'h0;
    1864: T381 = 1'h0;
    1865: T381 = 1'h0;
    1866: T381 = 1'h0;
    1867: T381 = 1'h0;
    1868: T381 = 1'h0;
    1869: T381 = 1'h0;
    1870: T381 = 1'h0;
    1871: T381 = 1'h0;
    1872: T381 = 1'h0;
    1873: T381 = 1'h0;
    1874: T381 = 1'h0;
    1875: T381 = 1'h0;
    1876: T381 = 1'h0;
    1877: T381 = 1'h0;
    1878: T381 = 1'h0;
    1879: T381 = 1'h0;
    1880: T381 = 1'h0;
    1881: T381 = 1'h0;
    1882: T381 = 1'h0;
    1883: T381 = 1'h0;
    1884: T381 = 1'h0;
    1885: T381 = 1'h0;
    1886: T381 = 1'h0;
    1887: T381 = 1'h0;
    1888: T381 = 1'h0;
    1889: T381 = 1'h0;
    1890: T381 = 1'h0;
    1891: T381 = 1'h0;
    1892: T381 = 1'h0;
    1893: T381 = 1'h0;
    1894: T381 = 1'h0;
    1895: T381 = 1'h0;
    1896: T381 = 1'h0;
    1897: T381 = 1'h0;
    1898: T381 = 1'h0;
    1899: T381 = 1'h0;
    1900: T381 = 1'h0;
    1901: T381 = 1'h0;
    1902: T381 = 1'h0;
    1903: T381 = 1'h0;
    1904: T381 = 1'h0;
    1905: T381 = 1'h0;
    1906: T381 = 1'h0;
    1907: T381 = 1'h0;
    1908: T381 = 1'h0;
    1909: T381 = 1'h0;
    1910: T381 = 1'h0;
    1911: T381 = 1'h0;
    1912: T381 = 1'h0;
    1913: T381 = 1'h0;
    1914: T381 = 1'h0;
    1915: T381 = 1'h0;
    1916: T381 = 1'h0;
    1917: T381 = 1'h0;
    1918: T381 = 1'h0;
    1919: T381 = 1'h0;
    1920: T381 = 1'h0;
    1921: T381 = 1'h0;
    1922: T381 = 1'h0;
    1923: T381 = 1'h0;
    1924: T381 = 1'h0;
    1925: T381 = 1'h0;
    1926: T381 = 1'h0;
    1927: T381 = 1'h0;
    1928: T381 = 1'h0;
    1929: T381 = 1'h0;
    1930: T381 = 1'h0;
    1931: T381 = 1'h0;
    1932: T381 = 1'h0;
    1933: T381 = 1'h0;
    1934: T381 = 1'h0;
    1935: T381 = 1'h0;
    1936: T381 = 1'h0;
    1937: T381 = 1'h0;
    1938: T381 = 1'h0;
    1939: T381 = 1'h0;
    1940: T381 = 1'h0;
    1941: T381 = 1'h0;
    1942: T381 = 1'h0;
    1943: T381 = 1'h0;
    1944: T381 = 1'h0;
    1945: T381 = 1'h0;
    1946: T381 = 1'h0;
    1947: T381 = 1'h0;
    1948: T381 = 1'h0;
    1949: T381 = 1'h0;
    1950: T381 = 1'h0;
    1951: T381 = 1'h0;
    1952: T381 = 1'h0;
    1953: T381 = 1'h0;
    1954: T381 = 1'h0;
    1955: T381 = 1'h0;
    1956: T381 = 1'h0;
    1957: T381 = 1'h0;
    1958: T381 = 1'h0;
    1959: T381 = 1'h0;
    1960: T381 = 1'h0;
    1961: T381 = 1'h0;
    1962: T381 = 1'h0;
    1963: T381 = 1'h0;
    1964: T381 = 1'h0;
    1965: T381 = 1'h0;
    1966: T381 = 1'h0;
    1967: T381 = 1'h0;
    1968: T381 = 1'h0;
    1969: T381 = 1'h0;
    1970: T381 = 1'h0;
    1971: T381 = 1'h0;
    1972: T381 = 1'h0;
    1973: T381 = 1'h0;
    1974: T381 = 1'h0;
    1975: T381 = 1'h0;
    1976: T381 = 1'h0;
    1977: T381 = 1'h0;
    1978: T381 = 1'h0;
    1979: T381 = 1'h0;
    1980: T381 = 1'h0;
    1981: T381 = 1'h0;
    1982: T381 = 1'h0;
    1983: T381 = 1'h0;
    1984: T381 = 1'h0;
    1985: T381 = 1'h0;
    1986: T381 = 1'h0;
    1987: T381 = 1'h0;
    1988: T381 = 1'h0;
    1989: T381 = 1'h0;
    1990: T381 = 1'h0;
    1991: T381 = 1'h0;
    1992: T381 = 1'h0;
    1993: T381 = 1'h0;
    1994: T381 = 1'h0;
    1995: T381 = 1'h0;
    1996: T381 = 1'h0;
    1997: T381 = 1'h0;
    1998: T381 = 1'h0;
    1999: T381 = 1'h0;
    2000: T381 = 1'h0;
    2001: T381 = 1'h0;
    2002: T381 = 1'h0;
    2003: T381 = 1'h0;
    2004: T381 = 1'h0;
    2005: T381 = 1'h0;
    2006: T381 = 1'h0;
    2007: T381 = 1'h0;
    2008: T381 = 1'h0;
    2009: T381 = 1'h0;
    2010: T381 = 1'h0;
    2011: T381 = 1'h0;
    2012: T381 = 1'h0;
    2013: T381 = 1'h0;
    2014: T381 = 1'h0;
    2015: T381 = 1'h0;
    2016: T381 = 1'h0;
    2017: T381 = 1'h0;
    2018: T381 = 1'h0;
    2019: T381 = 1'h0;
    2020: T381 = 1'h0;
    2021: T381 = 1'h0;
    2022: T381 = 1'h0;
    2023: T381 = 1'h0;
    2024: T381 = 1'h0;
    2025: T381 = 1'h0;
    2026: T381 = 1'h0;
    2027: T381 = 1'h0;
    2028: T381 = 1'h0;
    2029: T381 = 1'h0;
    2030: T381 = 1'h0;
    2031: T381 = 1'h0;
    2032: T381 = 1'h0;
    2033: T381 = 1'h0;
    2034: T381 = 1'h0;
    2035: T381 = 1'h0;
    2036: T381 = 1'h0;
    2037: T381 = 1'h0;
    2038: T381 = 1'h0;
    2039: T381 = 1'h0;
    2040: T381 = 1'h0;
    2041: T381 = 1'h0;
    2042: T381 = 1'h0;
    2043: T381 = 1'h0;
    2044: T381 = 1'h0;
    2045: T381 = 1'h0;
    2046: T381 = 1'h0;
    2047: T381 = 1'h0;
    2048: T381 = 1'h0;
    2049: T381 = 1'h0;
    2050: T381 = 1'h0;
    2051: T381 = 1'h0;
    2052: T381 = 1'h0;
    2053: T381 = 1'h0;
    2054: T381 = 1'h0;
    2055: T381 = 1'h0;
    2056: T381 = 1'h0;
    2057: T381 = 1'h0;
    2058: T381 = 1'h0;
    2059: T381 = 1'h0;
    2060: T381 = 1'h0;
    2061: T381 = 1'h0;
    2062: T381 = 1'h0;
    2063: T381 = 1'h0;
    2064: T381 = 1'h0;
    2065: T381 = 1'h0;
    2066: T381 = 1'h0;
    2067: T381 = 1'h0;
    2068: T381 = 1'h0;
    2069: T381 = 1'h0;
    2070: T381 = 1'h0;
    2071: T381 = 1'h0;
    2072: T381 = 1'h0;
    2073: T381 = 1'h0;
    2074: T381 = 1'h0;
    2075: T381 = 1'h0;
    2076: T381 = 1'h0;
    2077: T381 = 1'h0;
    2078: T381 = 1'h0;
    2079: T381 = 1'h0;
    2080: T381 = 1'h0;
    2081: T381 = 1'h0;
    2082: T381 = 1'h0;
    2083: T381 = 1'h0;
    2084: T381 = 1'h0;
    2085: T381 = 1'h0;
    2086: T381 = 1'h0;
    2087: T381 = 1'h0;
    2088: T381 = 1'h0;
    2089: T381 = 1'h0;
    2090: T381 = 1'h0;
    2091: T381 = 1'h0;
    2092: T381 = 1'h0;
    2093: T381 = 1'h0;
    2094: T381 = 1'h0;
    2095: T381 = 1'h0;
    2096: T381 = 1'h0;
    2097: T381 = 1'h0;
    2098: T381 = 1'h0;
    2099: T381 = 1'h0;
    2100: T381 = 1'h0;
    2101: T381 = 1'h0;
    2102: T381 = 1'h0;
    2103: T381 = 1'h0;
    2104: T381 = 1'h0;
    2105: T381 = 1'h0;
    2106: T381 = 1'h0;
    2107: T381 = 1'h0;
    2108: T381 = 1'h0;
    2109: T381 = 1'h0;
    2110: T381 = 1'h0;
    2111: T381 = 1'h0;
    2112: T381 = 1'h0;
    2113: T381 = 1'h0;
    2114: T381 = 1'h0;
    2115: T381 = 1'h0;
    2116: T381 = 1'h0;
    2117: T381 = 1'h0;
    2118: T381 = 1'h0;
    2119: T381 = 1'h0;
    2120: T381 = 1'h0;
    2121: T381 = 1'h0;
    2122: T381 = 1'h0;
    2123: T381 = 1'h0;
    2124: T381 = 1'h0;
    2125: T381 = 1'h0;
    2126: T381 = 1'h0;
    2127: T381 = 1'h0;
    2128: T381 = 1'h0;
    2129: T381 = 1'h0;
    2130: T381 = 1'h0;
    2131: T381 = 1'h0;
    2132: T381 = 1'h0;
    2133: T381 = 1'h0;
    2134: T381 = 1'h0;
    2135: T381 = 1'h0;
    2136: T381 = 1'h0;
    2137: T381 = 1'h0;
    2138: T381 = 1'h0;
    2139: T381 = 1'h0;
    2140: T381 = 1'h0;
    2141: T381 = 1'h0;
    2142: T381 = 1'h0;
    2143: T381 = 1'h0;
    2144: T381 = 1'h0;
    2145: T381 = 1'h0;
    2146: T381 = 1'h0;
    2147: T381 = 1'h0;
    2148: T381 = 1'h0;
    2149: T381 = 1'h0;
    2150: T381 = 1'h0;
    2151: T381 = 1'h0;
    2152: T381 = 1'h0;
    2153: T381 = 1'h0;
    2154: T381 = 1'h0;
    2155: T381 = 1'h0;
    2156: T381 = 1'h0;
    2157: T381 = 1'h0;
    2158: T381 = 1'h0;
    2159: T381 = 1'h0;
    2160: T381 = 1'h0;
    2161: T381 = 1'h0;
    2162: T381 = 1'h0;
    2163: T381 = 1'h0;
    2164: T381 = 1'h0;
    2165: T381 = 1'h0;
    2166: T381 = 1'h0;
    2167: T381 = 1'h0;
    2168: T381 = 1'h0;
    2169: T381 = 1'h0;
    2170: T381 = 1'h0;
    2171: T381 = 1'h0;
    2172: T381 = 1'h0;
    2173: T381 = 1'h0;
    2174: T381 = 1'h0;
    2175: T381 = 1'h0;
    2176: T381 = 1'h0;
    2177: T381 = 1'h0;
    2178: T381 = 1'h0;
    2179: T381 = 1'h0;
    2180: T381 = 1'h0;
    2181: T381 = 1'h0;
    2182: T381 = 1'h0;
    2183: T381 = 1'h0;
    2184: T381 = 1'h0;
    2185: T381 = 1'h0;
    2186: T381 = 1'h0;
    2187: T381 = 1'h0;
    2188: T381 = 1'h0;
    2189: T381 = 1'h0;
    2190: T381 = 1'h0;
    2191: T381 = 1'h0;
    2192: T381 = 1'h0;
    2193: T381 = 1'h0;
    2194: T381 = 1'h0;
    2195: T381 = 1'h0;
    2196: T381 = 1'h0;
    2197: T381 = 1'h0;
    2198: T381 = 1'h0;
    2199: T381 = 1'h0;
    2200: T381 = 1'h0;
    2201: T381 = 1'h0;
    2202: T381 = 1'h0;
    2203: T381 = 1'h0;
    2204: T381 = 1'h0;
    2205: T381 = 1'h0;
    2206: T381 = 1'h0;
    2207: T381 = 1'h0;
    2208: T381 = 1'h0;
    2209: T381 = 1'h0;
    2210: T381 = 1'h0;
    2211: T381 = 1'h0;
    2212: T381 = 1'h0;
    2213: T381 = 1'h0;
    2214: T381 = 1'h0;
    2215: T381 = 1'h0;
    2216: T381 = 1'h0;
    2217: T381 = 1'h0;
    2218: T381 = 1'h0;
    2219: T381 = 1'h0;
    2220: T381 = 1'h0;
    2221: T381 = 1'h0;
    2222: T381 = 1'h0;
    2223: T381 = 1'h0;
    2224: T381 = 1'h0;
    2225: T381 = 1'h0;
    2226: T381 = 1'h0;
    2227: T381 = 1'h0;
    2228: T381 = 1'h0;
    2229: T381 = 1'h0;
    2230: T381 = 1'h0;
    2231: T381 = 1'h0;
    2232: T381 = 1'h0;
    2233: T381 = 1'h0;
    2234: T381 = 1'h0;
    2235: T381 = 1'h0;
    2236: T381 = 1'h0;
    2237: T381 = 1'h0;
    2238: T381 = 1'h0;
    2239: T381 = 1'h0;
    2240: T381 = 1'h0;
    2241: T381 = 1'h0;
    2242: T381 = 1'h0;
    2243: T381 = 1'h0;
    2244: T381 = 1'h0;
    2245: T381 = 1'h0;
    2246: T381 = 1'h0;
    2247: T381 = 1'h0;
    2248: T381 = 1'h0;
    2249: T381 = 1'h0;
    2250: T381 = 1'h0;
    2251: T381 = 1'h0;
    2252: T381 = 1'h0;
    2253: T381 = 1'h0;
    2254: T381 = 1'h0;
    2255: T381 = 1'h0;
    2256: T381 = 1'h0;
    2257: T381 = 1'h0;
    2258: T381 = 1'h0;
    2259: T381 = 1'h0;
    2260: T381 = 1'h0;
    2261: T381 = 1'h0;
    2262: T381 = 1'h0;
    2263: T381 = 1'h0;
    2264: T381 = 1'h0;
    2265: T381 = 1'h0;
    2266: T381 = 1'h0;
    2267: T381 = 1'h0;
    2268: T381 = 1'h0;
    2269: T381 = 1'h0;
    2270: T381 = 1'h0;
    2271: T381 = 1'h0;
    2272: T381 = 1'h0;
    2273: T381 = 1'h0;
    2274: T381 = 1'h0;
    2275: T381 = 1'h0;
    2276: T381 = 1'h0;
    2277: T381 = 1'h0;
    2278: T381 = 1'h0;
    2279: T381 = 1'h0;
    2280: T381 = 1'h0;
    2281: T381 = 1'h0;
    2282: T381 = 1'h0;
    2283: T381 = 1'h0;
    2284: T381 = 1'h0;
    2285: T381 = 1'h0;
    2286: T381 = 1'h0;
    2287: T381 = 1'h0;
    2288: T381 = 1'h0;
    2289: T381 = 1'h0;
    2290: T381 = 1'h0;
    2291: T381 = 1'h0;
    2292: T381 = 1'h0;
    2293: T381 = 1'h0;
    2294: T381 = 1'h0;
    2295: T381 = 1'h0;
    2296: T381 = 1'h0;
    2297: T381 = 1'h0;
    2298: T381 = 1'h0;
    2299: T381 = 1'h0;
    2300: T381 = 1'h0;
    2301: T381 = 1'h0;
    2302: T381 = 1'h0;
    2303: T381 = 1'h0;
    2304: T381 = 1'h0;
    2305: T381 = 1'h0;
    2306: T381 = 1'h0;
    2307: T381 = 1'h0;
    2308: T381 = 1'h0;
    2309: T381 = 1'h0;
    2310: T381 = 1'h0;
    2311: T381 = 1'h0;
    2312: T381 = 1'h0;
    2313: T381 = 1'h0;
    2314: T381 = 1'h0;
    2315: T381 = 1'h0;
    2316: T381 = 1'h0;
    2317: T381 = 1'h0;
    2318: T381 = 1'h0;
    2319: T381 = 1'h0;
    2320: T381 = 1'h0;
    2321: T381 = 1'h0;
    2322: T381 = 1'h0;
    2323: T381 = 1'h0;
    2324: T381 = 1'h0;
    2325: T381 = 1'h0;
    2326: T381 = 1'h0;
    2327: T381 = 1'h0;
    2328: T381 = 1'h0;
    2329: T381 = 1'h0;
    2330: T381 = 1'h0;
    2331: T381 = 1'h0;
    2332: T381 = 1'h0;
    2333: T381 = 1'h0;
    2334: T381 = 1'h0;
    2335: T381 = 1'h0;
    2336: T381 = 1'h0;
    2337: T381 = 1'h0;
    2338: T381 = 1'h0;
    2339: T381 = 1'h0;
    2340: T381 = 1'h0;
    2341: T381 = 1'h0;
    2342: T381 = 1'h0;
    2343: T381 = 1'h0;
    2344: T381 = 1'h0;
    2345: T381 = 1'h0;
    2346: T381 = 1'h0;
    2347: T381 = 1'h0;
    2348: T381 = 1'h0;
    2349: T381 = 1'h0;
    2350: T381 = 1'h0;
    2351: T381 = 1'h0;
    2352: T381 = 1'h0;
    2353: T381 = 1'h0;
    2354: T381 = 1'h0;
    2355: T381 = 1'h0;
    2356: T381 = 1'h0;
    2357: T381 = 1'h0;
    2358: T381 = 1'h0;
    2359: T381 = 1'h0;
    2360: T381 = 1'h0;
    2361: T381 = 1'h0;
    2362: T381 = 1'h0;
    2363: T381 = 1'h0;
    2364: T381 = 1'h0;
    2365: T381 = 1'h0;
    2366: T381 = 1'h0;
    2367: T381 = 1'h0;
    2368: T381 = 1'h0;
    2369: T381 = 1'h0;
    2370: T381 = 1'h0;
    2371: T381 = 1'h0;
    2372: T381 = 1'h0;
    2373: T381 = 1'h0;
    2374: T381 = 1'h0;
    2375: T381 = 1'h0;
    2376: T381 = 1'h0;
    2377: T381 = 1'h0;
    2378: T381 = 1'h0;
    2379: T381 = 1'h0;
    2380: T381 = 1'h0;
    2381: T381 = 1'h0;
    2382: T381 = 1'h0;
    2383: T381 = 1'h0;
    2384: T381 = 1'h0;
    2385: T381 = 1'h0;
    2386: T381 = 1'h0;
    2387: T381 = 1'h0;
    2388: T381 = 1'h0;
    2389: T381 = 1'h0;
    2390: T381 = 1'h0;
    2391: T381 = 1'h0;
    2392: T381 = 1'h0;
    2393: T381 = 1'h0;
    2394: T381 = 1'h0;
    2395: T381 = 1'h0;
    2396: T381 = 1'h0;
    2397: T381 = 1'h0;
    2398: T381 = 1'h0;
    2399: T381 = 1'h0;
    2400: T381 = 1'h0;
    2401: T381 = 1'h0;
    2402: T381 = 1'h0;
    2403: T381 = 1'h0;
    2404: T381 = 1'h0;
    2405: T381 = 1'h0;
    2406: T381 = 1'h0;
    2407: T381 = 1'h0;
    2408: T381 = 1'h0;
    2409: T381 = 1'h0;
    2410: T381 = 1'h0;
    2411: T381 = 1'h0;
    2412: T381 = 1'h0;
    2413: T381 = 1'h0;
    2414: T381 = 1'h0;
    2415: T381 = 1'h0;
    2416: T381 = 1'h0;
    2417: T381 = 1'h0;
    2418: T381 = 1'h0;
    2419: T381 = 1'h0;
    2420: T381 = 1'h0;
    2421: T381 = 1'h0;
    2422: T381 = 1'h0;
    2423: T381 = 1'h0;
    2424: T381 = 1'h0;
    2425: T381 = 1'h0;
    2426: T381 = 1'h0;
    2427: T381 = 1'h0;
    2428: T381 = 1'h0;
    2429: T381 = 1'h0;
    2430: T381 = 1'h0;
    2431: T381 = 1'h0;
    2432: T381 = 1'h0;
    2433: T381 = 1'h0;
    2434: T381 = 1'h0;
    2435: T381 = 1'h0;
    2436: T381 = 1'h0;
    2437: T381 = 1'h0;
    2438: T381 = 1'h0;
    2439: T381 = 1'h0;
    2440: T381 = 1'h0;
    2441: T381 = 1'h0;
    2442: T381 = 1'h0;
    2443: T381 = 1'h0;
    2444: T381 = 1'h0;
    2445: T381 = 1'h0;
    2446: T381 = 1'h0;
    2447: T381 = 1'h0;
    2448: T381 = 1'h0;
    2449: T381 = 1'h0;
    2450: T381 = 1'h0;
    2451: T381 = 1'h0;
    2452: T381 = 1'h0;
    2453: T381 = 1'h0;
    2454: T381 = 1'h0;
    2455: T381 = 1'h0;
    2456: T381 = 1'h0;
    2457: T381 = 1'h0;
    2458: T381 = 1'h0;
    2459: T381 = 1'h0;
    2460: T381 = 1'h0;
    2461: T381 = 1'h0;
    2462: T381 = 1'h0;
    2463: T381 = 1'h0;
    2464: T381 = 1'h0;
    2465: T381 = 1'h0;
    2466: T381 = 1'h0;
    2467: T381 = 1'h0;
    2468: T381 = 1'h0;
    2469: T381 = 1'h0;
    2470: T381 = 1'h0;
    2471: T381 = 1'h0;
    2472: T381 = 1'h0;
    2473: T381 = 1'h0;
    2474: T381 = 1'h0;
    2475: T381 = 1'h0;
    2476: T381 = 1'h0;
    2477: T381 = 1'h0;
    2478: T381 = 1'h0;
    2479: T381 = 1'h0;
    2480: T381 = 1'h0;
    2481: T381 = 1'h0;
    2482: T381 = 1'h0;
    2483: T381 = 1'h0;
    2484: T381 = 1'h0;
    2485: T381 = 1'h0;
    2486: T381 = 1'h0;
    2487: T381 = 1'h0;
    2488: T381 = 1'h0;
    2489: T381 = 1'h0;
    2490: T381 = 1'h0;
    2491: T381 = 1'h0;
    2492: T381 = 1'h0;
    2493: T381 = 1'h0;
    2494: T381 = 1'h0;
    2495: T381 = 1'h0;
    2496: T381 = 1'h0;
    2497: T381 = 1'h0;
    2498: T381 = 1'h0;
    2499: T381 = 1'h0;
    2500: T381 = 1'h0;
    2501: T381 = 1'h0;
    2502: T381 = 1'h0;
    2503: T381 = 1'h0;
    2504: T381 = 1'h0;
    2505: T381 = 1'h0;
    2506: T381 = 1'h0;
    2507: T381 = 1'h0;
    2508: T381 = 1'h0;
    2509: T381 = 1'h0;
    2510: T381 = 1'h0;
    2511: T381 = 1'h0;
    2512: T381 = 1'h0;
    2513: T381 = 1'h0;
    2514: T381 = 1'h0;
    2515: T381 = 1'h0;
    2516: T381 = 1'h0;
    2517: T381 = 1'h0;
    2518: T381 = 1'h0;
    2519: T381 = 1'h0;
    2520: T381 = 1'h0;
    2521: T381 = 1'h0;
    2522: T381 = 1'h0;
    2523: T381 = 1'h0;
    2524: T381 = 1'h0;
    2525: T381 = 1'h0;
    2526: T381 = 1'h0;
    2527: T381 = 1'h0;
    2528: T381 = 1'h0;
    2529: T381 = 1'h0;
    2530: T381 = 1'h0;
    2531: T381 = 1'h0;
    2532: T381 = 1'h0;
    2533: T381 = 1'h0;
    2534: T381 = 1'h0;
    2535: T381 = 1'h0;
    2536: T381 = 1'h0;
    2537: T381 = 1'h0;
    2538: T381 = 1'h0;
    2539: T381 = 1'h0;
    2540: T381 = 1'h0;
    2541: T381 = 1'h0;
    2542: T381 = 1'h0;
    2543: T381 = 1'h0;
    2544: T381 = 1'h0;
    2545: T381 = 1'h0;
    2546: T381 = 1'h0;
    2547: T381 = 1'h0;
    2548: T381 = 1'h0;
    2549: T381 = 1'h0;
    2550: T381 = 1'h0;
    2551: T381 = 1'h0;
    2552: T381 = 1'h0;
    2553: T381 = 1'h0;
    2554: T381 = 1'h0;
    2555: T381 = 1'h0;
    2556: T381 = 1'h0;
    2557: T381 = 1'h0;
    2558: T381 = 1'h0;
    2559: T381 = 1'h0;
    2560: T381 = 1'h0;
    2561: T381 = 1'h0;
    2562: T381 = 1'h0;
    2563: T381 = 1'h0;
    2564: T381 = 1'h0;
    2565: T381 = 1'h0;
    2566: T381 = 1'h0;
    2567: T381 = 1'h0;
    2568: T381 = 1'h0;
    2569: T381 = 1'h0;
    2570: T381 = 1'h0;
    2571: T381 = 1'h0;
    2572: T381 = 1'h0;
    2573: T381 = 1'h0;
    2574: T381 = 1'h0;
    2575: T381 = 1'h0;
    2576: T381 = 1'h0;
    2577: T381 = 1'h0;
    2578: T381 = 1'h0;
    2579: T381 = 1'h0;
    2580: T381 = 1'h0;
    2581: T381 = 1'h0;
    2582: T381 = 1'h0;
    2583: T381 = 1'h0;
    2584: T381 = 1'h0;
    2585: T381 = 1'h0;
    2586: T381 = 1'h0;
    2587: T381 = 1'h0;
    2588: T381 = 1'h0;
    2589: T381 = 1'h0;
    2590: T381 = 1'h0;
    2591: T381 = 1'h0;
    2592: T381 = 1'h0;
    2593: T381 = 1'h0;
    2594: T381 = 1'h0;
    2595: T381 = 1'h0;
    2596: T381 = 1'h0;
    2597: T381 = 1'h0;
    2598: T381 = 1'h0;
    2599: T381 = 1'h0;
    2600: T381 = 1'h0;
    2601: T381 = 1'h0;
    2602: T381 = 1'h0;
    2603: T381 = 1'h0;
    2604: T381 = 1'h0;
    2605: T381 = 1'h0;
    2606: T381 = 1'h0;
    2607: T381 = 1'h0;
    2608: T381 = 1'h0;
    2609: T381 = 1'h0;
    2610: T381 = 1'h0;
    2611: T381 = 1'h0;
    2612: T381 = 1'h0;
    2613: T381 = 1'h0;
    2614: T381 = 1'h0;
    2615: T381 = 1'h0;
    2616: T381 = 1'h0;
    2617: T381 = 1'h0;
    2618: T381 = 1'h0;
    2619: T381 = 1'h0;
    2620: T381 = 1'h0;
    2621: T381 = 1'h0;
    2622: T381 = 1'h0;
    2623: T381 = 1'h0;
    2624: T381 = 1'h0;
    2625: T381 = 1'h0;
    2626: T381 = 1'h0;
    2627: T381 = 1'h0;
    2628: T381 = 1'h0;
    2629: T381 = 1'h0;
    2630: T381 = 1'h0;
    2631: T381 = 1'h0;
    2632: T381 = 1'h0;
    2633: T381 = 1'h0;
    2634: T381 = 1'h0;
    2635: T381 = 1'h0;
    2636: T381 = 1'h0;
    2637: T381 = 1'h0;
    2638: T381 = 1'h0;
    2639: T381 = 1'h0;
    2640: T381 = 1'h0;
    2641: T381 = 1'h0;
    2642: T381 = 1'h0;
    2643: T381 = 1'h0;
    2644: T381 = 1'h0;
    2645: T381 = 1'h0;
    2646: T381 = 1'h0;
    2647: T381 = 1'h0;
    2648: T381 = 1'h0;
    2649: T381 = 1'h0;
    2650: T381 = 1'h0;
    2651: T381 = 1'h0;
    2652: T381 = 1'h0;
    2653: T381 = 1'h0;
    2654: T381 = 1'h0;
    2655: T381 = 1'h0;
    2656: T381 = 1'h0;
    2657: T381 = 1'h0;
    2658: T381 = 1'h0;
    2659: T381 = 1'h0;
    2660: T381 = 1'h0;
    2661: T381 = 1'h0;
    2662: T381 = 1'h0;
    2663: T381 = 1'h0;
    2664: T381 = 1'h0;
    2665: T381 = 1'h0;
    2666: T381 = 1'h0;
    2667: T381 = 1'h0;
    2668: T381 = 1'h0;
    2669: T381 = 1'h0;
    2670: T381 = 1'h0;
    2671: T381 = 1'h0;
    2672: T381 = 1'h0;
    2673: T381 = 1'h0;
    2674: T381 = 1'h0;
    2675: T381 = 1'h0;
    2676: T381 = 1'h0;
    2677: T381 = 1'h0;
    2678: T381 = 1'h0;
    2679: T381 = 1'h0;
    2680: T381 = 1'h0;
    2681: T381 = 1'h0;
    2682: T381 = 1'h0;
    2683: T381 = 1'h0;
    2684: T381 = 1'h0;
    2685: T381 = 1'h0;
    2686: T381 = 1'h0;
    2687: T381 = 1'h0;
    2688: T381 = 1'h0;
    2689: T381 = 1'h0;
    2690: T381 = 1'h0;
    2691: T381 = 1'h0;
    2692: T381 = 1'h0;
    2693: T381 = 1'h0;
    2694: T381 = 1'h0;
    2695: T381 = 1'h0;
    2696: T381 = 1'h0;
    2697: T381 = 1'h0;
    2698: T381 = 1'h0;
    2699: T381 = 1'h0;
    2700: T381 = 1'h0;
    2701: T381 = 1'h0;
    2702: T381 = 1'h0;
    2703: T381 = 1'h0;
    2704: T381 = 1'h0;
    2705: T381 = 1'h0;
    2706: T381 = 1'h0;
    2707: T381 = 1'h0;
    2708: T381 = 1'h0;
    2709: T381 = 1'h0;
    2710: T381 = 1'h0;
    2711: T381 = 1'h0;
    2712: T381 = 1'h0;
    2713: T381 = 1'h0;
    2714: T381 = 1'h0;
    2715: T381 = 1'h0;
    2716: T381 = 1'h0;
    2717: T381 = 1'h0;
    2718: T381 = 1'h0;
    2719: T381 = 1'h0;
    2720: T381 = 1'h0;
    2721: T381 = 1'h0;
    2722: T381 = 1'h0;
    2723: T381 = 1'h0;
    2724: T381 = 1'h0;
    2725: T381 = 1'h0;
    2726: T381 = 1'h0;
    2727: T381 = 1'h0;
    2728: T381 = 1'h0;
    2729: T381 = 1'h0;
    2730: T381 = 1'h0;
    2731: T381 = 1'h0;
    2732: T381 = 1'h0;
    2733: T381 = 1'h0;
    2734: T381 = 1'h0;
    2735: T381 = 1'h0;
    2736: T381 = 1'h0;
    2737: T381 = 1'h0;
    2738: T381 = 1'h0;
    2739: T381 = 1'h0;
    2740: T381 = 1'h0;
    2741: T381 = 1'h0;
    2742: T381 = 1'h0;
    2743: T381 = 1'h0;
    2744: T381 = 1'h0;
    2745: T381 = 1'h0;
    2746: T381 = 1'h0;
    2747: T381 = 1'h0;
    2748: T381 = 1'h0;
    2749: T381 = 1'h0;
    2750: T381 = 1'h0;
    2751: T381 = 1'h0;
    2752: T381 = 1'h0;
    2753: T381 = 1'h0;
    2754: T381 = 1'h0;
    2755: T381 = 1'h0;
    2756: T381 = 1'h0;
    2757: T381 = 1'h0;
    2758: T381 = 1'h0;
    2759: T381 = 1'h0;
    2760: T381 = 1'h0;
    2761: T381 = 1'h0;
    2762: T381 = 1'h0;
    2763: T381 = 1'h0;
    2764: T381 = 1'h0;
    2765: T381 = 1'h0;
    2766: T381 = 1'h0;
    2767: T381 = 1'h0;
    2768: T381 = 1'h0;
    2769: T381 = 1'h0;
    2770: T381 = 1'h0;
    2771: T381 = 1'h0;
    2772: T381 = 1'h0;
    2773: T381 = 1'h0;
    2774: T381 = 1'h0;
    2775: T381 = 1'h0;
    2776: T381 = 1'h0;
    2777: T381 = 1'h0;
    2778: T381 = 1'h0;
    2779: T381 = 1'h0;
    2780: T381 = 1'h0;
    2781: T381 = 1'h0;
    2782: T381 = 1'h0;
    2783: T381 = 1'h0;
    2784: T381 = 1'h0;
    2785: T381 = 1'h0;
    2786: T381 = 1'h0;
    2787: T381 = 1'h0;
    2788: T381 = 1'h0;
    2789: T381 = 1'h0;
    2790: T381 = 1'h0;
    2791: T381 = 1'h0;
    2792: T381 = 1'h0;
    2793: T381 = 1'h0;
    2794: T381 = 1'h0;
    2795: T381 = 1'h0;
    2796: T381 = 1'h0;
    2797: T381 = 1'h0;
    2798: T381 = 1'h0;
    2799: T381 = 1'h0;
    2800: T381 = 1'h0;
    2801: T381 = 1'h0;
    2802: T381 = 1'h0;
    2803: T381 = 1'h0;
    2804: T381 = 1'h0;
    2805: T381 = 1'h0;
    2806: T381 = 1'h0;
    2807: T381 = 1'h0;
    2808: T381 = 1'h0;
    2809: T381 = 1'h0;
    2810: T381 = 1'h0;
    2811: T381 = 1'h0;
    2812: T381 = 1'h0;
    2813: T381 = 1'h0;
    2814: T381 = 1'h0;
    2815: T381 = 1'h0;
    2816: T381 = 1'h0;
    2817: T381 = 1'h0;
    2818: T381 = 1'h0;
    2819: T381 = 1'h0;
    2820: T381 = 1'h0;
    2821: T381 = 1'h0;
    2822: T381 = 1'h0;
    2823: T381 = 1'h0;
    2824: T381 = 1'h0;
    2825: T381 = 1'h0;
    2826: T381 = 1'h0;
    2827: T381 = 1'h0;
    2828: T381 = 1'h0;
    2829: T381 = 1'h0;
    2830: T381 = 1'h0;
    2831: T381 = 1'h0;
    2832: T381 = 1'h0;
    2833: T381 = 1'h0;
    2834: T381 = 1'h0;
    2835: T381 = 1'h0;
    2836: T381 = 1'h0;
    2837: T381 = 1'h0;
    2838: T381 = 1'h0;
    2839: T381 = 1'h0;
    2840: T381 = 1'h0;
    2841: T381 = 1'h0;
    2842: T381 = 1'h0;
    2843: T381 = 1'h0;
    2844: T381 = 1'h0;
    2845: T381 = 1'h0;
    2846: T381 = 1'h0;
    2847: T381 = 1'h0;
    2848: T381 = 1'h0;
    2849: T381 = 1'h0;
    2850: T381 = 1'h0;
    2851: T381 = 1'h0;
    2852: T381 = 1'h0;
    2853: T381 = 1'h0;
    2854: T381 = 1'h0;
    2855: T381 = 1'h0;
    2856: T381 = 1'h0;
    2857: T381 = 1'h0;
    2858: T381 = 1'h0;
    2859: T381 = 1'h0;
    2860: T381 = 1'h0;
    2861: T381 = 1'h0;
    2862: T381 = 1'h0;
    2863: T381 = 1'h0;
    2864: T381 = 1'h0;
    2865: T381 = 1'h0;
    2866: T381 = 1'h0;
    2867: T381 = 1'h0;
    2868: T381 = 1'h0;
    2869: T381 = 1'h0;
    2870: T381 = 1'h0;
    2871: T381 = 1'h0;
    2872: T381 = 1'h0;
    2873: T381 = 1'h0;
    2874: T381 = 1'h0;
    2875: T381 = 1'h0;
    2876: T381 = 1'h0;
    2877: T381 = 1'h0;
    2878: T381 = 1'h0;
    2879: T381 = 1'h0;
    2880: T381 = 1'h0;
    2881: T381 = 1'h0;
    2882: T381 = 1'h0;
    2883: T381 = 1'h0;
    2884: T381 = 1'h0;
    2885: T381 = 1'h0;
    2886: T381 = 1'h0;
    2887: T381 = 1'h0;
    2888: T381 = 1'h0;
    2889: T381 = 1'h0;
    2890: T381 = 1'h0;
    2891: T381 = 1'h0;
    2892: T381 = 1'h0;
    2893: T381 = 1'h0;
    2894: T381 = 1'h0;
    2895: T381 = 1'h0;
    2896: T381 = 1'h0;
    2897: T381 = 1'h0;
    2898: T381 = 1'h0;
    2899: T381 = 1'h0;
    2900: T381 = 1'h0;
    2901: T381 = 1'h0;
    2902: T381 = 1'h0;
    2903: T381 = 1'h0;
    2904: T381 = 1'h0;
    2905: T381 = 1'h0;
    2906: T381 = 1'h0;
    2907: T381 = 1'h0;
    2908: T381 = 1'h0;
    2909: T381 = 1'h0;
    2910: T381 = 1'h0;
    2911: T381 = 1'h0;
    2912: T381 = 1'h0;
    2913: T381 = 1'h0;
    2914: T381 = 1'h0;
    2915: T381 = 1'h0;
    2916: T381 = 1'h0;
    2917: T381 = 1'h0;
    2918: T381 = 1'h0;
    2919: T381 = 1'h0;
    2920: T381 = 1'h0;
    2921: T381 = 1'h0;
    2922: T381 = 1'h0;
    2923: T381 = 1'h0;
    2924: T381 = 1'h0;
    2925: T381 = 1'h0;
    2926: T381 = 1'h0;
    2927: T381 = 1'h0;
    2928: T381 = 1'h0;
    2929: T381 = 1'h0;
    2930: T381 = 1'h0;
    2931: T381 = 1'h0;
    2932: T381 = 1'h0;
    2933: T381 = 1'h0;
    2934: T381 = 1'h0;
    2935: T381 = 1'h0;
    2936: T381 = 1'h0;
    2937: T381 = 1'h0;
    2938: T381 = 1'h0;
    2939: T381 = 1'h0;
    2940: T381 = 1'h0;
    2941: T381 = 1'h0;
    2942: T381 = 1'h0;
    2943: T381 = 1'h0;
    2944: T381 = 1'h0;
    2945: T381 = 1'h0;
    2946: T381 = 1'h0;
    2947: T381 = 1'h0;
    2948: T381 = 1'h0;
    2949: T381 = 1'h0;
    2950: T381 = 1'h0;
    2951: T381 = 1'h0;
    2952: T381 = 1'h0;
    2953: T381 = 1'h0;
    2954: T381 = 1'h0;
    2955: T381 = 1'h0;
    2956: T381 = 1'h0;
    2957: T381 = 1'h0;
    2958: T381 = 1'h0;
    2959: T381 = 1'h0;
    2960: T381 = 1'h0;
    2961: T381 = 1'h0;
    2962: T381 = 1'h0;
    2963: T381 = 1'h0;
    2964: T381 = 1'h0;
    2965: T381 = 1'h0;
    2966: T381 = 1'h0;
    2967: T381 = 1'h0;
    2968: T381 = 1'h0;
    2969: T381 = 1'h0;
    2970: T381 = 1'h0;
    2971: T381 = 1'h0;
    2972: T381 = 1'h0;
    2973: T381 = 1'h0;
    2974: T381 = 1'h0;
    2975: T381 = 1'h0;
    2976: T381 = 1'h0;
    2977: T381 = 1'h0;
    2978: T381 = 1'h0;
    2979: T381 = 1'h0;
    2980: T381 = 1'h0;
    2981: T381 = 1'h0;
    2982: T381 = 1'h0;
    2983: T381 = 1'h0;
    2984: T381 = 1'h0;
    2985: T381 = 1'h0;
    2986: T381 = 1'h0;
    2987: T381 = 1'h0;
    2988: T381 = 1'h0;
    2989: T381 = 1'h0;
    2990: T381 = 1'h0;
    2991: T381 = 1'h0;
    2992: T381 = 1'h0;
    2993: T381 = 1'h0;
    2994: T381 = 1'h0;
    2995: T381 = 1'h0;
    2996: T381 = 1'h0;
    2997: T381 = 1'h0;
    2998: T381 = 1'h0;
    2999: T381 = 1'h0;
    3000: T381 = 1'h0;
    3001: T381 = 1'h0;
    3002: T381 = 1'h0;
    3003: T381 = 1'h0;
    3004: T381 = 1'h0;
    3005: T381 = 1'h0;
    3006: T381 = 1'h0;
    3007: T381 = 1'h0;
    3008: T381 = 1'h0;
    3009: T381 = 1'h0;
    3010: T381 = 1'h0;
    3011: T381 = 1'h0;
    3012: T381 = 1'h0;
    3013: T381 = 1'h0;
    3014: T381 = 1'h0;
    3015: T381 = 1'h0;
    3016: T381 = 1'h0;
    3017: T381 = 1'h0;
    3018: T381 = 1'h0;
    3019: T381 = 1'h0;
    3020: T381 = 1'h0;
    3021: T381 = 1'h0;
    3022: T381 = 1'h0;
    3023: T381 = 1'h0;
    3024: T381 = 1'h0;
    3025: T381 = 1'h0;
    3026: T381 = 1'h0;
    3027: T381 = 1'h0;
    3028: T381 = 1'h0;
    3029: T381 = 1'h0;
    3030: T381 = 1'h0;
    3031: T381 = 1'h0;
    3032: T381 = 1'h0;
    3033: T381 = 1'h0;
    3034: T381 = 1'h0;
    3035: T381 = 1'h0;
    3036: T381 = 1'h0;
    3037: T381 = 1'h0;
    3038: T381 = 1'h0;
    3039: T381 = 1'h0;
    3040: T381 = 1'h0;
    3041: T381 = 1'h0;
    3042: T381 = 1'h0;
    3043: T381 = 1'h0;
    3044: T381 = 1'h0;
    3045: T381 = 1'h0;
    3046: T381 = 1'h0;
    3047: T381 = 1'h0;
    3048: T381 = 1'h0;
    3049: T381 = 1'h0;
    3050: T381 = 1'h0;
    3051: T381 = 1'h0;
    3052: T381 = 1'h0;
    3053: T381 = 1'h0;
    3054: T381 = 1'h0;
    3055: T381 = 1'h0;
    3056: T381 = 1'h0;
    3057: T381 = 1'h0;
    3058: T381 = 1'h0;
    3059: T381 = 1'h0;
    3060: T381 = 1'h0;
    3061: T381 = 1'h0;
    3062: T381 = 1'h0;
    3063: T381 = 1'h0;
    3064: T381 = 1'h0;
    3065: T381 = 1'h0;
    3066: T381 = 1'h0;
    3067: T381 = 1'h0;
    3068: T381 = 1'h0;
    3069: T381 = 1'h0;
    3070: T381 = 1'h0;
    3071: T381 = 1'h0;
    3072: T381 = 1'h1;
    3073: T381 = 1'h1;
    3074: T381 = 1'h1;
    3075: T381 = 1'h0;
    3076: T381 = 1'h0;
    3077: T381 = 1'h0;
    3078: T381 = 1'h0;
    3079: T381 = 1'h0;
    3080: T381 = 1'h0;
    3081: T381 = 1'h0;
    3082: T381 = 1'h0;
    3083: T381 = 1'h0;
    3084: T381 = 1'h0;
    3085: T381 = 1'h0;
    3086: T381 = 1'h0;
    3087: T381 = 1'h0;
    3088: T381 = 1'h0;
    3089: T381 = 1'h0;
    3090: T381 = 1'h0;
    3091: T381 = 1'h0;
    3092: T381 = 1'h0;
    3093: T381 = 1'h0;
    3094: T381 = 1'h0;
    3095: T381 = 1'h0;
    3096: T381 = 1'h0;
    3097: T381 = 1'h0;
    3098: T381 = 1'h0;
    3099: T381 = 1'h0;
    3100: T381 = 1'h0;
    3101: T381 = 1'h0;
    3102: T381 = 1'h0;
    3103: T381 = 1'h0;
    3104: T381 = 1'h0;
    3105: T381 = 1'h0;
    3106: T381 = 1'h0;
    3107: T381 = 1'h0;
    3108: T381 = 1'h0;
    3109: T381 = 1'h0;
    3110: T381 = 1'h0;
    3111: T381 = 1'h0;
    3112: T381 = 1'h0;
    3113: T381 = 1'h0;
    3114: T381 = 1'h0;
    3115: T381 = 1'h0;
    3116: T381 = 1'h0;
    3117: T381 = 1'h0;
    3118: T381 = 1'h0;
    3119: T381 = 1'h0;
    3120: T381 = 1'h0;
    3121: T381 = 1'h0;
    3122: T381 = 1'h0;
    3123: T381 = 1'h0;
    3124: T381 = 1'h0;
    3125: T381 = 1'h0;
    3126: T381 = 1'h0;
    3127: T381 = 1'h0;
    3128: T381 = 1'h0;
    3129: T381 = 1'h0;
    3130: T381 = 1'h0;
    3131: T381 = 1'h0;
    3132: T381 = 1'h0;
    3133: T381 = 1'h0;
    3134: T381 = 1'h0;
    3135: T381 = 1'h0;
    3136: T381 = 1'h0;
    3137: T381 = 1'h0;
    3138: T381 = 1'h0;
    3139: T381 = 1'h0;
    3140: T381 = 1'h0;
    3141: T381 = 1'h0;
    3142: T381 = 1'h0;
    3143: T381 = 1'h0;
    3144: T381 = 1'h0;
    3145: T381 = 1'h0;
    3146: T381 = 1'h0;
    3147: T381 = 1'h0;
    3148: T381 = 1'h0;
    3149: T381 = 1'h0;
    3150: T381 = 1'h0;
    3151: T381 = 1'h0;
    3152: T381 = 1'h0;
    3153: T381 = 1'h0;
    3154: T381 = 1'h0;
    3155: T381 = 1'h0;
    3156: T381 = 1'h0;
    3157: T381 = 1'h0;
    3158: T381 = 1'h0;
    3159: T381 = 1'h0;
    3160: T381 = 1'h0;
    3161: T381 = 1'h0;
    3162: T381 = 1'h0;
    3163: T381 = 1'h0;
    3164: T381 = 1'h0;
    3165: T381 = 1'h0;
    3166: T381 = 1'h0;
    3167: T381 = 1'h0;
    3168: T381 = 1'h0;
    3169: T381 = 1'h0;
    3170: T381 = 1'h0;
    3171: T381 = 1'h0;
    3172: T381 = 1'h0;
    3173: T381 = 1'h0;
    3174: T381 = 1'h0;
    3175: T381 = 1'h0;
    3176: T381 = 1'h0;
    3177: T381 = 1'h0;
    3178: T381 = 1'h0;
    3179: T381 = 1'h0;
    3180: T381 = 1'h0;
    3181: T381 = 1'h0;
    3182: T381 = 1'h0;
    3183: T381 = 1'h0;
    3184: T381 = 1'h0;
    3185: T381 = 1'h0;
    3186: T381 = 1'h0;
    3187: T381 = 1'h0;
    3188: T381 = 1'h0;
    3189: T381 = 1'h0;
    3190: T381 = 1'h0;
    3191: T381 = 1'h0;
    3192: T381 = 1'h0;
    3193: T381 = 1'h0;
    3194: T381 = 1'h0;
    3195: T381 = 1'h0;
    3196: T381 = 1'h0;
    3197: T381 = 1'h0;
    3198: T381 = 1'h0;
    3199: T381 = 1'h0;
    3200: T381 = 1'h0;
    3201: T381 = 1'h0;
    3202: T381 = 1'h0;
    3203: T381 = 1'h0;
    3204: T381 = 1'h0;
    3205: T381 = 1'h0;
    3206: T381 = 1'h0;
    3207: T381 = 1'h0;
    3208: T381 = 1'h0;
    3209: T381 = 1'h0;
    3210: T381 = 1'h0;
    3211: T381 = 1'h0;
    3212: T381 = 1'h0;
    3213: T381 = 1'h0;
    3214: T381 = 1'h0;
    3215: T381 = 1'h0;
    3216: T381 = 1'h0;
    3217: T381 = 1'h0;
    3218: T381 = 1'h0;
    3219: T381 = 1'h0;
    3220: T381 = 1'h0;
    3221: T381 = 1'h0;
    3222: T381 = 1'h0;
    3223: T381 = 1'h0;
    3224: T381 = 1'h0;
    3225: T381 = 1'h0;
    3226: T381 = 1'h0;
    3227: T381 = 1'h0;
    3228: T381 = 1'h0;
    3229: T381 = 1'h0;
    3230: T381 = 1'h0;
    3231: T381 = 1'h0;
    3232: T381 = 1'h0;
    3233: T381 = 1'h0;
    3234: T381 = 1'h0;
    3235: T381 = 1'h0;
    3236: T381 = 1'h0;
    3237: T381 = 1'h0;
    3238: T381 = 1'h0;
    3239: T381 = 1'h0;
    3240: T381 = 1'h0;
    3241: T381 = 1'h0;
    3242: T381 = 1'h0;
    3243: T381 = 1'h0;
    3244: T381 = 1'h0;
    3245: T381 = 1'h0;
    3246: T381 = 1'h0;
    3247: T381 = 1'h0;
    3248: T381 = 1'h0;
    3249: T381 = 1'h0;
    3250: T381 = 1'h0;
    3251: T381 = 1'h0;
    3252: T381 = 1'h0;
    3253: T381 = 1'h0;
    3254: T381 = 1'h0;
    3255: T381 = 1'h0;
    3256: T381 = 1'h0;
    3257: T381 = 1'h0;
    3258: T381 = 1'h0;
    3259: T381 = 1'h0;
    3260: T381 = 1'h0;
    3261: T381 = 1'h0;
    3262: T381 = 1'h0;
    3263: T381 = 1'h0;
    3264: T381 = 1'h1;
    3265: T381 = 1'h1;
    3266: T381 = 1'h1;
    3267: T381 = 1'h1;
    3268: T381 = 1'h1;
    3269: T381 = 1'h1;
    3270: T381 = 1'h1;
    3271: T381 = 1'h1;
    3272: T381 = 1'h1;
    3273: T381 = 1'h1;
    3274: T381 = 1'h1;
    3275: T381 = 1'h1;
    3276: T381 = 1'h1;
    3277: T381 = 1'h1;
    3278: T381 = 1'h1;
    3279: T381 = 1'h1;
    3280: T381 = 1'h0;
    3281: T381 = 1'h0;
    3282: T381 = 1'h0;
    3283: T381 = 1'h0;
    3284: T381 = 1'h0;
    3285: T381 = 1'h0;
    3286: T381 = 1'h0;
    3287: T381 = 1'h0;
    3288: T381 = 1'h0;
    3289: T381 = 1'h0;
    3290: T381 = 1'h0;
    3291: T381 = 1'h0;
    3292: T381 = 1'h0;
    3293: T381 = 1'h0;
    3294: T381 = 1'h0;
    3295: T381 = 1'h0;
    3296: T381 = 1'h0;
    3297: T381 = 1'h0;
    3298: T381 = 1'h0;
    3299: T381 = 1'h0;
    3300: T381 = 1'h0;
    3301: T381 = 1'h0;
    3302: T381 = 1'h0;
    3303: T381 = 1'h0;
    3304: T381 = 1'h0;
    3305: T381 = 1'h0;
    3306: T381 = 1'h0;
    3307: T381 = 1'h0;
    3308: T381 = 1'h0;
    3309: T381 = 1'h0;
    3310: T381 = 1'h0;
    3311: T381 = 1'h0;
    3312: T381 = 1'h0;
    3313: T381 = 1'h0;
    3314: T381 = 1'h0;
    3315: T381 = 1'h0;
    3316: T381 = 1'h0;
    3317: T381 = 1'h0;
    3318: T381 = 1'h0;
    3319: T381 = 1'h0;
    3320: T381 = 1'h0;
    3321: T381 = 1'h0;
    3322: T381 = 1'h0;
    3323: T381 = 1'h0;
    3324: T381 = 1'h0;
    3325: T381 = 1'h0;
    3326: T381 = 1'h0;
    3327: T381 = 1'h0;
    3328: T381 = 1'h0;
    3329: T381 = 1'h0;
    3330: T381 = 1'h0;
    3331: T381 = 1'h0;
    3332: T381 = 1'h0;
    3333: T381 = 1'h0;
    3334: T381 = 1'h0;
    3335: T381 = 1'h0;
    3336: T381 = 1'h0;
    3337: T381 = 1'h0;
    3338: T381 = 1'h0;
    3339: T381 = 1'h0;
    3340: T381 = 1'h0;
    3341: T381 = 1'h0;
    3342: T381 = 1'h0;
    3343: T381 = 1'h0;
    3344: T381 = 1'h0;
    3345: T381 = 1'h0;
    3346: T381 = 1'h0;
    3347: T381 = 1'h0;
    3348: T381 = 1'h0;
    3349: T381 = 1'h0;
    3350: T381 = 1'h0;
    3351: T381 = 1'h0;
    3352: T381 = 1'h0;
    3353: T381 = 1'h0;
    3354: T381 = 1'h0;
    3355: T381 = 1'h0;
    3356: T381 = 1'h0;
    3357: T381 = 1'h0;
    3358: T381 = 1'h0;
    3359: T381 = 1'h0;
    3360: T381 = 1'h0;
    3361: T381 = 1'h0;
    3362: T381 = 1'h0;
    3363: T381 = 1'h0;
    3364: T381 = 1'h0;
    3365: T381 = 1'h0;
    3366: T381 = 1'h0;
    3367: T381 = 1'h0;
    3368: T381 = 1'h0;
    3369: T381 = 1'h0;
    3370: T381 = 1'h0;
    3371: T381 = 1'h0;
    3372: T381 = 1'h0;
    3373: T381 = 1'h0;
    3374: T381 = 1'h0;
    3375: T381 = 1'h0;
    3376: T381 = 1'h0;
    3377: T381 = 1'h0;
    3378: T381 = 1'h0;
    3379: T381 = 1'h0;
    3380: T381 = 1'h0;
    3381: T381 = 1'h0;
    3382: T381 = 1'h0;
    3383: T381 = 1'h0;
    3384: T381 = 1'h0;
    3385: T381 = 1'h0;
    3386: T381 = 1'h0;
    3387: T381 = 1'h0;
    3388: T381 = 1'h0;
    3389: T381 = 1'h0;
    3390: T381 = 1'h0;
    3391: T381 = 1'h0;
    3392: T381 = 1'h0;
    3393: T381 = 1'h0;
    3394: T381 = 1'h0;
    3395: T381 = 1'h0;
    3396: T381 = 1'h0;
    3397: T381 = 1'h0;
    3398: T381 = 1'h0;
    3399: T381 = 1'h0;
    3400: T381 = 1'h0;
    3401: T381 = 1'h0;
    3402: T381 = 1'h0;
    3403: T381 = 1'h0;
    3404: T381 = 1'h0;
    3405: T381 = 1'h0;
    3406: T381 = 1'h0;
    3407: T381 = 1'h0;
    3408: T381 = 1'h0;
    3409: T381 = 1'h0;
    3410: T381 = 1'h0;
    3411: T381 = 1'h0;
    3412: T381 = 1'h0;
    3413: T381 = 1'h0;
    3414: T381 = 1'h0;
    3415: T381 = 1'h0;
    3416: T381 = 1'h0;
    3417: T381 = 1'h0;
    3418: T381 = 1'h0;
    3419: T381 = 1'h0;
    3420: T381 = 1'h0;
    3421: T381 = 1'h0;
    3422: T381 = 1'h0;
    3423: T381 = 1'h0;
    3424: T381 = 1'h0;
    3425: T381 = 1'h0;
    3426: T381 = 1'h0;
    3427: T381 = 1'h0;
    3428: T381 = 1'h0;
    3429: T381 = 1'h0;
    3430: T381 = 1'h0;
    3431: T381 = 1'h0;
    3432: T381 = 1'h0;
    3433: T381 = 1'h0;
    3434: T381 = 1'h0;
    3435: T381 = 1'h0;
    3436: T381 = 1'h0;
    3437: T381 = 1'h0;
    3438: T381 = 1'h0;
    3439: T381 = 1'h0;
    3440: T381 = 1'h0;
    3441: T381 = 1'h0;
    3442: T381 = 1'h0;
    3443: T381 = 1'h0;
    3444: T381 = 1'h0;
    3445: T381 = 1'h0;
    3446: T381 = 1'h0;
    3447: T381 = 1'h0;
    3448: T381 = 1'h0;
    3449: T381 = 1'h0;
    3450: T381 = 1'h0;
    3451: T381 = 1'h0;
    3452: T381 = 1'h0;
    3453: T381 = 1'h0;
    3454: T381 = 1'h0;
    3455: T381 = 1'h0;
    3456: T381 = 1'h0;
    3457: T381 = 1'h0;
    3458: T381 = 1'h0;
    3459: T381 = 1'h0;
    3460: T381 = 1'h0;
    3461: T381 = 1'h0;
    3462: T381 = 1'h0;
    3463: T381 = 1'h0;
    3464: T381 = 1'h0;
    3465: T381 = 1'h0;
    3466: T381 = 1'h0;
    3467: T381 = 1'h0;
    3468: T381 = 1'h0;
    3469: T381 = 1'h0;
    3470: T381 = 1'h0;
    3471: T381 = 1'h0;
    3472: T381 = 1'h0;
    3473: T381 = 1'h0;
    3474: T381 = 1'h0;
    3475: T381 = 1'h0;
    3476: T381 = 1'h0;
    3477: T381 = 1'h0;
    3478: T381 = 1'h0;
    3479: T381 = 1'h0;
    3480: T381 = 1'h0;
    3481: T381 = 1'h0;
    3482: T381 = 1'h0;
    3483: T381 = 1'h0;
    3484: T381 = 1'h0;
    3485: T381 = 1'h0;
    3486: T381 = 1'h0;
    3487: T381 = 1'h0;
    3488: T381 = 1'h0;
    3489: T381 = 1'h0;
    3490: T381 = 1'h0;
    3491: T381 = 1'h0;
    3492: T381 = 1'h0;
    3493: T381 = 1'h0;
    3494: T381 = 1'h0;
    3495: T381 = 1'h0;
    3496: T381 = 1'h0;
    3497: T381 = 1'h0;
    3498: T381 = 1'h0;
    3499: T381 = 1'h0;
    3500: T381 = 1'h0;
    3501: T381 = 1'h0;
    3502: T381 = 1'h0;
    3503: T381 = 1'h0;
    3504: T381 = 1'h0;
    3505: T381 = 1'h0;
    3506: T381 = 1'h0;
    3507: T381 = 1'h0;
    3508: T381 = 1'h0;
    3509: T381 = 1'h0;
    3510: T381 = 1'h0;
    3511: T381 = 1'h0;
    3512: T381 = 1'h0;
    3513: T381 = 1'h0;
    3514: T381 = 1'h0;
    3515: T381 = 1'h0;
    3516: T381 = 1'h0;
    3517: T381 = 1'h0;
    3518: T381 = 1'h0;
    3519: T381 = 1'h0;
    3520: T381 = 1'h0;
    3521: T381 = 1'h0;
    3522: T381 = 1'h0;
    3523: T381 = 1'h0;
    3524: T381 = 1'h0;
    3525: T381 = 1'h0;
    3526: T381 = 1'h0;
    3527: T381 = 1'h0;
    3528: T381 = 1'h0;
    3529: T381 = 1'h0;
    3530: T381 = 1'h0;
    3531: T381 = 1'h0;
    3532: T381 = 1'h0;
    3533: T381 = 1'h0;
    3534: T381 = 1'h0;
    3535: T381 = 1'h0;
    3536: T381 = 1'h0;
    3537: T381 = 1'h0;
    3538: T381 = 1'h0;
    3539: T381 = 1'h0;
    3540: T381 = 1'h0;
    3541: T381 = 1'h0;
    3542: T381 = 1'h0;
    3543: T381 = 1'h0;
    3544: T381 = 1'h0;
    3545: T381 = 1'h0;
    3546: T381 = 1'h0;
    3547: T381 = 1'h0;
    3548: T381 = 1'h0;
    3549: T381 = 1'h0;
    3550: T381 = 1'h0;
    3551: T381 = 1'h0;
    3552: T381 = 1'h0;
    3553: T381 = 1'h0;
    3554: T381 = 1'h0;
    3555: T381 = 1'h0;
    3556: T381 = 1'h0;
    3557: T381 = 1'h0;
    3558: T381 = 1'h0;
    3559: T381 = 1'h0;
    3560: T381 = 1'h0;
    3561: T381 = 1'h0;
    3562: T381 = 1'h0;
    3563: T381 = 1'h0;
    3564: T381 = 1'h0;
    3565: T381 = 1'h0;
    3566: T381 = 1'h0;
    3567: T381 = 1'h0;
    3568: T381 = 1'h0;
    3569: T381 = 1'h0;
    3570: T381 = 1'h0;
    3571: T381 = 1'h0;
    3572: T381 = 1'h0;
    3573: T381 = 1'h0;
    3574: T381 = 1'h0;
    3575: T381 = 1'h0;
    3576: T381 = 1'h0;
    3577: T381 = 1'h0;
    3578: T381 = 1'h0;
    3579: T381 = 1'h0;
    3580: T381 = 1'h0;
    3581: T381 = 1'h0;
    3582: T381 = 1'h0;
    3583: T381 = 1'h0;
    3584: T381 = 1'h0;
    3585: T381 = 1'h0;
    3586: T381 = 1'h0;
    3587: T381 = 1'h0;
    3588: T381 = 1'h0;
    3589: T381 = 1'h0;
    3590: T381 = 1'h0;
    3591: T381 = 1'h0;
    3592: T381 = 1'h0;
    3593: T381 = 1'h0;
    3594: T381 = 1'h0;
    3595: T381 = 1'h0;
    3596: T381 = 1'h0;
    3597: T381 = 1'h0;
    3598: T381 = 1'h0;
    3599: T381 = 1'h0;
    3600: T381 = 1'h0;
    3601: T381 = 1'h0;
    3602: T381 = 1'h0;
    3603: T381 = 1'h0;
    3604: T381 = 1'h0;
    3605: T381 = 1'h0;
    3606: T381 = 1'h0;
    3607: T381 = 1'h0;
    3608: T381 = 1'h0;
    3609: T381 = 1'h0;
    3610: T381 = 1'h0;
    3611: T381 = 1'h0;
    3612: T381 = 1'h0;
    3613: T381 = 1'h0;
    3614: T381 = 1'h0;
    3615: T381 = 1'h0;
    3616: T381 = 1'h0;
    3617: T381 = 1'h0;
    3618: T381 = 1'h0;
    3619: T381 = 1'h0;
    3620: T381 = 1'h0;
    3621: T381 = 1'h0;
    3622: T381 = 1'h0;
    3623: T381 = 1'h0;
    3624: T381 = 1'h0;
    3625: T381 = 1'h0;
    3626: T381 = 1'h0;
    3627: T381 = 1'h0;
    3628: T381 = 1'h0;
    3629: T381 = 1'h0;
    3630: T381 = 1'h0;
    3631: T381 = 1'h0;
    3632: T381 = 1'h0;
    3633: T381 = 1'h0;
    3634: T381 = 1'h0;
    3635: T381 = 1'h0;
    3636: T381 = 1'h0;
    3637: T381 = 1'h0;
    3638: T381 = 1'h0;
    3639: T381 = 1'h0;
    3640: T381 = 1'h0;
    3641: T381 = 1'h0;
    3642: T381 = 1'h0;
    3643: T381 = 1'h0;
    3644: T381 = 1'h0;
    3645: T381 = 1'h0;
    3646: T381 = 1'h0;
    3647: T381 = 1'h0;
    3648: T381 = 1'h0;
    3649: T381 = 1'h0;
    3650: T381 = 1'h0;
    3651: T381 = 1'h0;
    3652: T381 = 1'h0;
    3653: T381 = 1'h0;
    3654: T381 = 1'h0;
    3655: T381 = 1'h0;
    3656: T381 = 1'h0;
    3657: T381 = 1'h0;
    3658: T381 = 1'h0;
    3659: T381 = 1'h0;
    3660: T381 = 1'h0;
    3661: T381 = 1'h0;
    3662: T381 = 1'h0;
    3663: T381 = 1'h0;
    3664: T381 = 1'h0;
    3665: T381 = 1'h0;
    3666: T381 = 1'h0;
    3667: T381 = 1'h0;
    3668: T381 = 1'h0;
    3669: T381 = 1'h0;
    3670: T381 = 1'h0;
    3671: T381 = 1'h0;
    3672: T381 = 1'h0;
    3673: T381 = 1'h0;
    3674: T381 = 1'h0;
    3675: T381 = 1'h0;
    3676: T381 = 1'h0;
    3677: T381 = 1'h0;
    3678: T381 = 1'h0;
    3679: T381 = 1'h0;
    3680: T381 = 1'h0;
    3681: T381 = 1'h0;
    3682: T381 = 1'h0;
    3683: T381 = 1'h0;
    3684: T381 = 1'h0;
    3685: T381 = 1'h0;
    3686: T381 = 1'h0;
    3687: T381 = 1'h0;
    3688: T381 = 1'h0;
    3689: T381 = 1'h0;
    3690: T381 = 1'h0;
    3691: T381 = 1'h0;
    3692: T381 = 1'h0;
    3693: T381 = 1'h0;
    3694: T381 = 1'h0;
    3695: T381 = 1'h0;
    3696: T381 = 1'h0;
    3697: T381 = 1'h0;
    3698: T381 = 1'h0;
    3699: T381 = 1'h0;
    3700: T381 = 1'h0;
    3701: T381 = 1'h0;
    3702: T381 = 1'h0;
    3703: T381 = 1'h0;
    3704: T381 = 1'h0;
    3705: T381 = 1'h0;
    3706: T381 = 1'h0;
    3707: T381 = 1'h0;
    3708: T381 = 1'h0;
    3709: T381 = 1'h0;
    3710: T381 = 1'h0;
    3711: T381 = 1'h0;
    3712: T381 = 1'h0;
    3713: T381 = 1'h0;
    3714: T381 = 1'h0;
    3715: T381 = 1'h0;
    3716: T381 = 1'h0;
    3717: T381 = 1'h0;
    3718: T381 = 1'h0;
    3719: T381 = 1'h0;
    3720: T381 = 1'h0;
    3721: T381 = 1'h0;
    3722: T381 = 1'h0;
    3723: T381 = 1'h0;
    3724: T381 = 1'h0;
    3725: T381 = 1'h0;
    3726: T381 = 1'h0;
    3727: T381 = 1'h0;
    3728: T381 = 1'h0;
    3729: T381 = 1'h0;
    3730: T381 = 1'h0;
    3731: T381 = 1'h0;
    3732: T381 = 1'h0;
    3733: T381 = 1'h0;
    3734: T381 = 1'h0;
    3735: T381 = 1'h0;
    3736: T381 = 1'h0;
    3737: T381 = 1'h0;
    3738: T381 = 1'h0;
    3739: T381 = 1'h0;
    3740: T381 = 1'h0;
    3741: T381 = 1'h0;
    3742: T381 = 1'h0;
    3743: T381 = 1'h0;
    3744: T381 = 1'h0;
    3745: T381 = 1'h0;
    3746: T381 = 1'h0;
    3747: T381 = 1'h0;
    3748: T381 = 1'h0;
    3749: T381 = 1'h0;
    3750: T381 = 1'h0;
    3751: T381 = 1'h0;
    3752: T381 = 1'h0;
    3753: T381 = 1'h0;
    3754: T381 = 1'h0;
    3755: T381 = 1'h0;
    3756: T381 = 1'h0;
    3757: T381 = 1'h0;
    3758: T381 = 1'h0;
    3759: T381 = 1'h0;
    3760: T381 = 1'h0;
    3761: T381 = 1'h0;
    3762: T381 = 1'h0;
    3763: T381 = 1'h0;
    3764: T381 = 1'h0;
    3765: T381 = 1'h0;
    3766: T381 = 1'h0;
    3767: T381 = 1'h0;
    3768: T381 = 1'h0;
    3769: T381 = 1'h0;
    3770: T381 = 1'h0;
    3771: T381 = 1'h0;
    3772: T381 = 1'h0;
    3773: T381 = 1'h0;
    3774: T381 = 1'h0;
    3775: T381 = 1'h0;
    3776: T381 = 1'h0;
    3777: T381 = 1'h0;
    3778: T381 = 1'h0;
    3779: T381 = 1'h0;
    3780: T381 = 1'h0;
    3781: T381 = 1'h0;
    3782: T381 = 1'h0;
    3783: T381 = 1'h0;
    3784: T381 = 1'h0;
    3785: T381 = 1'h0;
    3786: T381 = 1'h0;
    3787: T381 = 1'h0;
    3788: T381 = 1'h0;
    3789: T381 = 1'h0;
    3790: T381 = 1'h0;
    3791: T381 = 1'h0;
    3792: T381 = 1'h0;
    3793: T381 = 1'h0;
    3794: T381 = 1'h0;
    3795: T381 = 1'h0;
    3796: T381 = 1'h0;
    3797: T381 = 1'h0;
    3798: T381 = 1'h0;
    3799: T381 = 1'h0;
    3800: T381 = 1'h0;
    3801: T381 = 1'h0;
    3802: T381 = 1'h0;
    3803: T381 = 1'h0;
    3804: T381 = 1'h0;
    3805: T381 = 1'h0;
    3806: T381 = 1'h0;
    3807: T381 = 1'h0;
    3808: T381 = 1'h0;
    3809: T381 = 1'h0;
    3810: T381 = 1'h0;
    3811: T381 = 1'h0;
    3812: T381 = 1'h0;
    3813: T381 = 1'h0;
    3814: T381 = 1'h0;
    3815: T381 = 1'h0;
    3816: T381 = 1'h0;
    3817: T381 = 1'h0;
    3818: T381 = 1'h0;
    3819: T381 = 1'h0;
    3820: T381 = 1'h0;
    3821: T381 = 1'h0;
    3822: T381 = 1'h0;
    3823: T381 = 1'h0;
    3824: T381 = 1'h0;
    3825: T381 = 1'h0;
    3826: T381 = 1'h0;
    3827: T381 = 1'h0;
    3828: T381 = 1'h0;
    3829: T381 = 1'h0;
    3830: T381 = 1'h0;
    3831: T381 = 1'h0;
    3832: T381 = 1'h0;
    3833: T381 = 1'h0;
    3834: T381 = 1'h0;
    3835: T381 = 1'h0;
    3836: T381 = 1'h0;
    3837: T381 = 1'h0;
    3838: T381 = 1'h0;
    3839: T381 = 1'h0;
    3840: T381 = 1'h0;
    3841: T381 = 1'h0;
    3842: T381 = 1'h0;
    3843: T381 = 1'h0;
    3844: T381 = 1'h0;
    3845: T381 = 1'h0;
    3846: T381 = 1'h0;
    3847: T381 = 1'h0;
    3848: T381 = 1'h0;
    3849: T381 = 1'h0;
    3850: T381 = 1'h0;
    3851: T381 = 1'h0;
    3852: T381 = 1'h0;
    3853: T381 = 1'h0;
    3854: T381 = 1'h0;
    3855: T381 = 1'h0;
    3856: T381 = 1'h0;
    3857: T381 = 1'h0;
    3858: T381 = 1'h0;
    3859: T381 = 1'h0;
    3860: T381 = 1'h0;
    3861: T381 = 1'h0;
    3862: T381 = 1'h0;
    3863: T381 = 1'h0;
    3864: T381 = 1'h0;
    3865: T381 = 1'h0;
    3866: T381 = 1'h0;
    3867: T381 = 1'h0;
    3868: T381 = 1'h0;
    3869: T381 = 1'h0;
    3870: T381 = 1'h0;
    3871: T381 = 1'h0;
    3872: T381 = 1'h0;
    3873: T381 = 1'h0;
    3874: T381 = 1'h0;
    3875: T381 = 1'h0;
    3876: T381 = 1'h0;
    3877: T381 = 1'h0;
    3878: T381 = 1'h0;
    3879: T381 = 1'h0;
    3880: T381 = 1'h0;
    3881: T381 = 1'h0;
    3882: T381 = 1'h0;
    3883: T381 = 1'h0;
    3884: T381 = 1'h0;
    3885: T381 = 1'h0;
    3886: T381 = 1'h0;
    3887: T381 = 1'h0;
    3888: T381 = 1'h0;
    3889: T381 = 1'h0;
    3890: T381 = 1'h0;
    3891: T381 = 1'h0;
    3892: T381 = 1'h0;
    3893: T381 = 1'h0;
    3894: T381 = 1'h0;
    3895: T381 = 1'h0;
    3896: T381 = 1'h0;
    3897: T381 = 1'h0;
    3898: T381 = 1'h0;
    3899: T381 = 1'h0;
    3900: T381 = 1'h0;
    3901: T381 = 1'h0;
    3902: T381 = 1'h0;
    3903: T381 = 1'h0;
    3904: T381 = 1'h0;
    3905: T381 = 1'h0;
    3906: T381 = 1'h0;
    3907: T381 = 1'h0;
    3908: T381 = 1'h0;
    3909: T381 = 1'h0;
    3910: T381 = 1'h0;
    3911: T381 = 1'h0;
    3912: T381 = 1'h0;
    3913: T381 = 1'h0;
    3914: T381 = 1'h0;
    3915: T381 = 1'h0;
    3916: T381 = 1'h0;
    3917: T381 = 1'h0;
    3918: T381 = 1'h0;
    3919: T381 = 1'h0;
    3920: T381 = 1'h0;
    3921: T381 = 1'h0;
    3922: T381 = 1'h0;
    3923: T381 = 1'h0;
    3924: T381 = 1'h0;
    3925: T381 = 1'h0;
    3926: T381 = 1'h0;
    3927: T381 = 1'h0;
    3928: T381 = 1'h0;
    3929: T381 = 1'h0;
    3930: T381 = 1'h0;
    3931: T381 = 1'h0;
    3932: T381 = 1'h0;
    3933: T381 = 1'h0;
    3934: T381 = 1'h0;
    3935: T381 = 1'h0;
    3936: T381 = 1'h0;
    3937: T381 = 1'h0;
    3938: T381 = 1'h0;
    3939: T381 = 1'h0;
    3940: T381 = 1'h0;
    3941: T381 = 1'h0;
    3942: T381 = 1'h0;
    3943: T381 = 1'h0;
    3944: T381 = 1'h0;
    3945: T381 = 1'h0;
    3946: T381 = 1'h0;
    3947: T381 = 1'h0;
    3948: T381 = 1'h0;
    3949: T381 = 1'h0;
    3950: T381 = 1'h0;
    3951: T381 = 1'h0;
    3952: T381 = 1'h0;
    3953: T381 = 1'h0;
    3954: T381 = 1'h0;
    3955: T381 = 1'h0;
    3956: T381 = 1'h0;
    3957: T381 = 1'h0;
    3958: T381 = 1'h0;
    3959: T381 = 1'h0;
    3960: T381 = 1'h0;
    3961: T381 = 1'h0;
    3962: T381 = 1'h0;
    3963: T381 = 1'h0;
    3964: T381 = 1'h0;
    3965: T381 = 1'h0;
    3966: T381 = 1'h0;
    3967: T381 = 1'h0;
    3968: T381 = 1'h0;
    3969: T381 = 1'h0;
    3970: T381 = 1'h0;
    3971: T381 = 1'h0;
    3972: T381 = 1'h0;
    3973: T381 = 1'h0;
    3974: T381 = 1'h0;
    3975: T381 = 1'h0;
    3976: T381 = 1'h0;
    3977: T381 = 1'h0;
    3978: T381 = 1'h0;
    3979: T381 = 1'h0;
    3980: T381 = 1'h0;
    3981: T381 = 1'h0;
    3982: T381 = 1'h0;
    3983: T381 = 1'h0;
    3984: T381 = 1'h0;
    3985: T381 = 1'h0;
    3986: T381 = 1'h0;
    3987: T381 = 1'h0;
    3988: T381 = 1'h0;
    3989: T381 = 1'h0;
    3990: T381 = 1'h0;
    3991: T381 = 1'h0;
    3992: T381 = 1'h0;
    3993: T381 = 1'h0;
    3994: T381 = 1'h0;
    3995: T381 = 1'h0;
    3996: T381 = 1'h0;
    3997: T381 = 1'h0;
    3998: T381 = 1'h0;
    3999: T381 = 1'h0;
    4000: T381 = 1'h0;
    4001: T381 = 1'h0;
    4002: T381 = 1'h0;
    4003: T381 = 1'h0;
    4004: T381 = 1'h0;
    4005: T381 = 1'h0;
    4006: T381 = 1'h0;
    4007: T381 = 1'h0;
    4008: T381 = 1'h0;
    4009: T381 = 1'h0;
    4010: T381 = 1'h0;
    4011: T381 = 1'h0;
    4012: T381 = 1'h0;
    4013: T381 = 1'h0;
    4014: T381 = 1'h0;
    4015: T381 = 1'h0;
    4016: T381 = 1'h0;
    4017: T381 = 1'h0;
    4018: T381 = 1'h0;
    4019: T381 = 1'h0;
    4020: T381 = 1'h0;
    4021: T381 = 1'h0;
    4022: T381 = 1'h0;
    4023: T381 = 1'h0;
    4024: T381 = 1'h0;
    4025: T381 = 1'h0;
    4026: T381 = 1'h0;
    4027: T381 = 1'h0;
    4028: T381 = 1'h0;
    4029: T381 = 1'h0;
    4030: T381 = 1'h0;
    4031: T381 = 1'h0;
    4032: T381 = 1'h0;
    4033: T381 = 1'h0;
    4034: T381 = 1'h0;
    4035: T381 = 1'h0;
    4036: T381 = 1'h0;
    4037: T381 = 1'h0;
    4038: T381 = 1'h0;
    4039: T381 = 1'h0;
    4040: T381 = 1'h0;
    4041: T381 = 1'h0;
    4042: T381 = 1'h0;
    4043: T381 = 1'h0;
    4044: T381 = 1'h0;
    4045: T381 = 1'h0;
    4046: T381 = 1'h0;
    4047: T381 = 1'h0;
    4048: T381 = 1'h0;
    4049: T381 = 1'h0;
    4050: T381 = 1'h0;
    4051: T381 = 1'h0;
    4052: T381 = 1'h0;
    4053: T381 = 1'h0;
    4054: T381 = 1'h0;
    4055: T381 = 1'h0;
    4056: T381 = 1'h0;
    4057: T381 = 1'h0;
    4058: T381 = 1'h0;
    4059: T381 = 1'h0;
    4060: T381 = 1'h0;
    4061: T381 = 1'h0;
    4062: T381 = 1'h0;
    4063: T381 = 1'h0;
    4064: T381 = 1'h0;
    4065: T381 = 1'h0;
    4066: T381 = 1'h0;
    4067: T381 = 1'h0;
    4068: T381 = 1'h0;
    4069: T381 = 1'h0;
    4070: T381 = 1'h0;
    4071: T381 = 1'h0;
    4072: T381 = 1'h0;
    4073: T381 = 1'h0;
    4074: T381 = 1'h0;
    4075: T381 = 1'h0;
    4076: T381 = 1'h0;
    4077: T381 = 1'h0;
    4078: T381 = 1'h0;
    4079: T381 = 1'h0;
    4080: T381 = 1'h0;
    4081: T381 = 1'h0;
    4082: T381 = 1'h0;
    4083: T381 = 1'h0;
    4084: T381 = 1'h0;
    4085: T381 = 1'h0;
    4086: T381 = 1'h0;
    4087: T381 = 1'h0;
    4088: T381 = 1'h0;
    4089: T381 = 1'h0;
    4090: T381 = 1'h0;
    4091: T381 = 1'h0;
    4092: T381 = 1'h0;
    4093: T381 = 1'h0;
    4094: T381 = 1'h0;
    4095: T381 = 1'h0;
`ifndef SYNTHESIS
    default: T381 = {1{$random}};
`else
    default: T381 = 1'bx;
`endif
  endcase
  assign T383 = id_int_val ^ 1'h1;
  assign id_int_val = T386 | T384;
  assign T384 = T385 == 32'h33;
  assign T385 = io_dpath_inst & 32'hfc007077;
  assign T386 = T389 | T387;
  assign T387 = T388 == 32'h4063;
  assign T388 = io_dpath_inst & 32'h407f;
  assign T389 = T392 | T390;
  assign T390 = T391 == 32'h1063;
  assign T391 = io_dpath_inst & 32'h306f;
  assign T392 = T393 | T63;
  assign T393 = T394 | T66;
  assign T394 = T397 | T395;
  assign T395 = T396 == 32'h2004033;
  assign T396 = io_dpath_inst & 32'hfe004077;
  assign T397 = T400 | T398;
  assign T398 = T399 == 32'h5033;
  assign T399 = io_dpath_inst & 32'hbe007077;
  assign T400 = T403 | T401;
  assign T401 = T402 == 32'h501b;
  assign T402 = io_dpath_inst & 32'hbe00705f;
  assign T403 = T406 | T404;
  assign T404 = T405 == 32'h5013;
  assign T405 = io_dpath_inst & 32'hbc00707f;
  assign T406 = T409 | T407;
  assign T407 = T408 == 32'h2073;
  assign T408 = io_dpath_inst & 32'h207f;
  assign T409 = T410 | T69;
  assign T410 = T413 | T411;
  assign T411 = T412 == 32'h2013;
  assign T412 = io_dpath_inst & 32'h207f;
  assign T413 = T416 | T414;
  assign T414 = T415 == 32'h101b;
  assign T415 = io_dpath_inst & 32'hfe00305f;
  assign T416 = T419 | T417;
  assign T417 = T418 == 32'h1013;
  assign T418 = io_dpath_inst & 32'hfc00305f;
  assign T419 = T422 | T420;
  assign T420 = T421 == 32'h73;
  assign T421 = io_dpath_inst & 32'h7fffffff;
  assign T422 = T425 | T423;
  assign T423 = T424 == 32'h6f;
  assign T424 = io_dpath_inst & 32'h7f;
  assign T425 = T428 | T426;
  assign T426 = T427 == 32'h63;
  assign T427 = io_dpath_inst & 32'h707b;
  assign T428 = T431 | T429;
  assign T429 = T430 == 32'h33;
  assign T430 = io_dpath_inst & 32'hbe007077;
  assign T431 = T434 | T432;
  assign T432 = T433 == 32'h33;
  assign T433 = io_dpath_inst & 32'hfc00007f;
  assign T434 = T437 | T435;
  assign T435 = T436 == 32'h17;
  assign T436 = io_dpath_inst & 32'h5f;
  assign T437 = T440 | T438;
  assign T438 = T439 == 32'h13;
  assign T439 = io_dpath_inst & 32'h7077;
  assign T440 = T443 | T441;
  assign T441 = T442 == 32'hf;
  assign T442 = io_dpath_inst & 32'h607f;
  assign T443 = T446 | T444;
  assign T444 = T445 == 32'h3;
  assign T445 = io_dpath_inst & 32'h106f;
  assign T446 = T77 | T75;
  assign T447 = T448 | io_imem_resp_bits_xcpt_if;
  assign T448 = id_interrupt | io_imem_resp_bits_xcpt_ma;
  assign T449 = T450 & io_imem_resp_valid;
  assign T450 = id_interrupt & T451;
  assign T451 = take_pc ^ 1'h1;
  assign T452 = dcache_kill_mem | take_pc_wb;
  assign dcache_kill_mem = mem_reg_wen & io_dmem_replay_next_valid;
  assign T453 = replay_wb | wb_reg_xcpt;
  assign replay_wb = replay_wb_common | T454;
  assign T454 = wb_reg_rocc_val & T455;
  assign T455 = io_rocc_cmd_ready ^ 1'h1;
  assign replay_wb_common = T456 | io_dpath_csr_replay;
  assign T456 = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T457 = replay_mem & T458;
  assign T458 = take_pc_wb ^ 1'h1;
  assign replay_mem = T459 | fpu_kill_mem;
  assign T459 = dcache_kill_mem | mem_reg_replay;
  assign mem_xcpt = T461 | T460;
  assign T460 = mem_reg_mem_val & io_dmem_xcpt_pf_st;
  assign T461 = T463 | T462;
  assign T462 = mem_reg_mem_val & io_dmem_xcpt_pf_ld;
  assign T463 = T465 | T464;
  assign T464 = mem_reg_mem_val & io_dmem_xcpt_ma_st;
  assign T465 = T467 | T466;
  assign T466 = mem_reg_mem_val & io_dmem_xcpt_ma_ld;
  assign T467 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T468 = T470 & T469;
  assign T469 = mem_reg_replay_next ^ 1'h1;
  assign T470 = T471 & ex_reg_xcpt_interrupt;
  assign T471 = take_pc ^ 1'h1;
  assign io_rocc_s = io_dpath_status_s;
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign wb_rocc_val = wb_reg_rocc_val & T472;
  assign T472 = replay_wb_common ^ 1'h1;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = 1'h0;
  assign io_dmem_req_bits_cmd = ex_reg_mem_cmd;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_typ = ex_reg_mem_type;
  assign io_dmem_req_bits_kill = T473;
  assign T473 = killm_common | mem_xcpt;
  assign io_dmem_req_valid = ex_reg_mem_val;
  assign io_imem_invalidate = wb_reg_flush_inst;
  assign T474 = ctrl_killm ? 1'h0 : mem_reg_flush_inst;
  assign T475 = ctrl_killx ? 1'h0 : ex_reg_flush_inst;
  assign T476 = ctrl_killd ? 1'h0 : id_fence_i;
  assign io_imem_btb_update_bits_incorrectTarget = take_pc_mem;
  assign io_imem_btb_update_bits_isReturn = T477;
  assign T477 = mem_reg_jalr & io_dpath_mem_rs1_ra;
  assign io_imem_btb_update_bits_isCall = T478;
  assign T478 = mem_reg_wen & T479;
  assign T479 = io_dpath_mem_waddr[1'h0:1'h0];
  assign io_imem_btb_update_bits_isJump = T480;
  assign T480 = mem_reg_jal | mem_reg_jalr;
  assign io_imem_btb_update_bits_taken = T481;
  assign T481 = mem_reg_jal | T482;
  assign T482 = mem_reg_branch & io_dpath_mem_br_taken;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T483 = T486 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T484 = T485 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T485 = T246 & io_imem_btb_resp_valid;
  assign T486 = T278 & ex_reg_btb_hit;
  assign T487 = ctrl_killd ? 1'h0 : io_imem_btb_resp_valid;
  assign io_imem_btb_update_bits_prediction_bits_bht_index = mem_reg_btb_resp_bht_index;
  assign T488 = T486 ? ex_reg_btb_resp_bht_index : mem_reg_btb_resp_bht_index;
  assign T489 = T485 ? io_imem_btb_resp_bits_bht_index : ex_reg_btb_resp_bht_index;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T490 = T486 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T491 = T485 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T492 = T486 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T493 = T485 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T494 = T486 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T495 = T485 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T496 = T278 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T497;
  assign T497 = T498 | mem_reg_jalr;
  assign T498 = mem_reg_branch | mem_reg_jal;
  assign io_imem_resp_ready = T499;
  assign T499 = T500 | ctrl_draind;
  assign T500 = ctrl_stalld ^ 1'h1;
  assign io_imem_req_valid = take_pc;
  assign io_dpath_badvaddr_wen = wb_reg_xcpt;
  assign io_dpath_cause = wb_reg_cause;
  assign T501 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T467 ? mem_reg_cause : T667;
  assign T667 = {60'h0, T502};
  assign T502 = T466 ? 4'h8 : T503;
  assign T503 = T464 ? 4'h9 : T504;
  assign T504 = T462 ? 4'ha : 4'hb;
  assign T505 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T351 ? ex_reg_cause : 64'h2;
  assign T506 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = id_interrupt ? id_interrupt_cause : T668;
  assign T668 = {60'h0, T507};
  assign T507 = io_imem_resp_bits_xcpt_ma ? 4'h0 : T508;
  assign T508 = io_imem_resp_bits_xcpt_if ? 4'h1 : T509;
  assign T509 = T379 ? 4'h2 : T510;
  assign T510 = id_csr_privileged ? 4'h3 : T511;
  assign T511 = T355 ? 4'h3 : T512;
  assign T512 = id_syscall ? 4'h6 : 4'hc;
  assign id_interrupt_cause = T56 ? 64'h8000000000000000 : T513;
  assign T513 = T53 ? 64'h8000000000000001 : T514;
  assign T514 = T49 ? 64'h8000000000000002 : T515;
  assign T515 = T45 ? 64'h8000000000000003 : T516;
  assign T516 = T41 ? 64'h8000000000000004 : T517;
  assign T517 = T37 ? 64'h8000000000000005 : T518;
  assign T518 = T33 ? 64'h8000000000000006 : 64'h8000000000000007;
  assign io_dpath_exception = wb_reg_xcpt;
  assign io_dpath_retire = T519;
  assign T519 = wb_reg_valid & T520;
  assign T520 = replay_wb ^ 1'h1;
  assign T521 = ctrl_killm ? 1'h0 : mem_reg_valid;
  assign io_dpath_ll_ready = T522;
  assign T522 = wb_reg_wen ^ 1'h1;
  assign io_dpath_bypass_src_0 = T523;
  assign T523 = T532 ? 2'h0 : T524;
  assign T524 = T530 ? 2'h1 : T525;
  assign T525 = T526 ? 2'h2 : 2'h3;
  assign T526 = T528 & T527;
  assign T527 = io_dpath_mem_waddr == id_raddr1;
  assign T528 = mem_reg_wen & T529;
  assign T529 = mem_reg_mem_val ^ 1'h1;
  assign T530 = ex_reg_wen & T531;
  assign T531 = io_dpath_ex_waddr == id_raddr1;
  assign T532 = 5'h0 == id_raddr1;
  assign io_dpath_bypass_src_1 = T533;
  assign T533 = T540 ? 2'h0 : T534;
  assign T534 = T538 ? 2'h1 : T535;
  assign T535 = T536 ? 2'h2 : 2'h3;
  assign T536 = T528 & T537;
  assign T537 = io_dpath_mem_waddr == id_raddr2;
  assign T538 = ex_reg_wen & T539;
  assign T539 = io_dpath_ex_waddr == id_raddr2;
  assign T540 = 5'h0 == id_raddr2;
  assign io_dpath_bypass_0 = T541;
  assign T541 = T544 | T542;
  assign T542 = mem_reg_wen & T543;
  assign T543 = io_dpath_mem_waddr == id_raddr1;
  assign T544 = T545 | T526;
  assign T545 = T532 | T530;
  assign io_dpath_bypass_1 = T546;
  assign T546 = T549 | T547;
  assign T547 = mem_reg_wen & T548;
  assign T548 = io_dpath_mem_waddr == id_raddr2;
  assign T549 = T550 | T536;
  assign T550 = T540 | T538;
  assign io_dpath_mem_rocc_val = mem_reg_rocc_val;
  assign io_dpath_ex_rocc_val = ex_reg_rocc_val;
  assign io_dpath_ex_rs2_val = T551;
  assign T551 = T552 | ex_reg_rocc_val;
  assign T552 = ex_reg_mem_val & T553;
  assign T553 = T557 | T554;
  assign T554 = T556 | T555;
  assign T555 = ex_reg_mem_cmd == 5'h4;
  assign T556 = ex_reg_mem_cmd[2'h3:2'h3];
  assign T557 = T559 | T558;
  assign T558 = ex_reg_mem_cmd == 5'h7;
  assign T559 = ex_reg_mem_cmd == 5'h1;
  assign io_dpath_ex_mem_type = ex_reg_mem_type;
  assign io_dpath_wb_wen = T560;
  assign T560 = wb_reg_wen & T561;
  assign T561 = replay_wb ^ 1'h1;
  assign io_dpath_mem_wen = mem_reg_wen;
  assign io_dpath_mem_branch = mem_reg_branch;
  assign io_dpath_mem_jalr = mem_reg_jalr;
  assign io_dpath_ex_valid = ex_reg_valid;
  assign io_dpath_ex_wen = ex_reg_wen;
  assign io_dpath_mem_fp_val = mem_reg_fp_val;
  assign io_dpath_ex_fp_val = ex_reg_fp_val;
  assign io_dpath_wb_load = T562;
  assign T562 = wb_reg_mem_val & wb_reg_wen;
  assign io_dpath_mem_load = T563;
  assign T563 = mem_reg_mem_val & mem_reg_wen;
  assign io_dpath_sret = wb_reg_sret;
  assign io_dpath_csr = T669;
  assign T669 = {1'h0, wb_reg_csr};
  assign T564 = ctrl_killm ? 2'h0 : mem_reg_csr;
  assign io_dpath_div_mul_kill = T565;
  assign T565 = mem_reg_div_mul_val & killm_common;
  assign io_dpath_div_mul_val = ex_reg_div_mul_val;
  assign io_dpath_fn_alu = T566;
  assign T566 = id_fn_alu;
  assign id_fn_alu = {T602, T567};
  assign T567 = {T591, T568};
  assign T568 = {T577, T569};
  assign T569 = T572 | T570;
  assign T570 = T571 == 32'h7000;
  assign T571 = io_dpath_inst & 32'h7044;
  assign T572 = T575 | T573;
  assign T573 = T574 == 32'h1040;
  assign T574 = io_dpath_inst & 32'h1058;
  assign T575 = T576 == 32'h1010;
  assign T576 = io_dpath_inst & 32'h3054;
  assign T577 = T580 | T578;
  assign T578 = T579 == 32'h40001010;
  assign T579 = io_dpath_inst & 32'h40001054;
  assign T580 = T583 | T581;
  assign T581 = T582 == 32'h40000030;
  assign T582 = io_dpath_inst & 32'h40003034;
  assign T583 = T586 | T584;
  assign T584 = T585 == 32'h6010;
  assign T585 = io_dpath_inst & 32'h6054;
  assign T586 = T589 | T587;
  assign T587 = T588 == 32'h3010;
  assign T588 = io_dpath_inst & 32'h3054;
  assign T589 = T590 == 32'h2040;
  assign T590 = io_dpath_inst & 32'h2058;
  assign T591 = T594 | T592;
  assign T592 = T593 == 32'h4040;
  assign T593 = io_dpath_inst & 32'h4058;
  assign T594 = T597 | T595;
  assign T595 = T596 == 32'h4010;
  assign T596 = io_dpath_inst & 32'h5054;
  assign T597 = T600 | T598;
  assign T598 = T599 == 32'h4010;
  assign T599 = io_dpath_inst & 32'h40004054;
  assign T600 = T601 == 32'h2010;
  assign T601 = io_dpath_inst & 32'h2054;
  assign T602 = T605 | T603;
  assign T603 = T604 == 32'h40001010;
  assign T604 = io_dpath_inst & 32'h40003054;
  assign T605 = T606 | T581;
  assign T606 = id_branch | T607;
  assign T607 = T608 == 32'h2010;
  assign T608 = io_dpath_inst & 32'h6054;
  assign io_dpath_fn_dw = T609;
  assign T609 = id_fn_dw;
  assign id_fn_dw = T612 | T610;
  assign T610 = T611 == 32'h0;
  assign T611 = io_dpath_inst & 32'h8;
  assign T612 = T613 == 32'h0;
  assign T613 = io_dpath_inst & 32'h10;
  assign io_dpath_sel_imm = T614;
  assign T614 = id_sel_imm;
  assign id_sel_imm = {T624, T615};
  assign T615 = {T621, T616};
  assign T616 = T619 | T617;
  assign T617 = T618 == 32'h40;
  assign T618 = io_dpath_inst & 32'h44;
  assign T619 = T620 == 32'h8;
  assign T620 = io_dpath_inst & 32'h18;
  assign T621 = T622 | T619;
  assign T622 = T623 == 32'h4;
  assign T623 = io_dpath_inst & 32'h44;
  assign T624 = T627 | T625;
  assign T625 = T626 == 32'h10;
  assign T626 = io_dpath_inst & 32'h14;
  assign T627 = T628 | id_jalr;
  assign T628 = T629 == 32'h0;
  assign T629 = io_dpath_inst & 32'h24;
  assign io_dpath_sel_alu1 = T630;
  assign T630 = id_sel_alu1;
  assign id_sel_alu1 = {T638, T631};
  assign T631 = T632 | T179;
  assign T632 = T633 | T181;
  assign T633 = T636 | T634;
  assign T634 = T635 == 32'h0;
  assign T635 = io_dpath_inst & 32'h50;
  assign T636 = T637 == 32'h0;
  assign T637 = io_dpath_inst & 32'h4004;
  assign T638 = T639 | id_jal;
  assign T639 = T640 == 32'h4;
  assign T640 = io_dpath_inst & 32'h24;
  assign io_dpath_sel_alu2 = T670;
  assign T670 = {1'h0, T641};
  assign T641 = id_sel_alu2;
  assign id_sel_alu2 = {T652, T642};
  assign T642 = T645 | T643;
  assign T643 = T644 == 32'h4050;
  assign T644 = io_dpath_inst & 32'h4050;
  assign T645 = T646 | id_jal;
  assign T646 = T647 | T144;
  assign T647 = T650 | T648;
  assign T648 = T649 == 32'h0;
  assign T649 = io_dpath_inst & 32'h20;
  assign T650 = T651 == 32'h0;
  assign T651 = io_dpath_inst & 32'h58;
  assign T652 = T655 | T653;
  assign T653 = T654 == 32'h4000;
  assign T654 = io_dpath_inst & 32'h4008;
  assign T655 = T656 | T179;
  assign T656 = T657 | T181;
  assign T657 = T658 == 32'h0;
  assign T658 = io_dpath_inst & 32'h48;
  assign io_dpath_ren_0 = id_renx1;
  assign io_dpath_ren_1 = id_renx2;
  assign io_dpath_killd = T659;
  assign T659 = take_pc | T660;
  assign T660 = ctrl_stalld & T661;
  assign T661 = ctrl_draind ^ 1'h1;
  assign io_dpath_sel_pc = T671;
  assign T671 = {1'h0, T662};
  assign T662 = wb_reg_xcpt ? 2'h3 : T663;
  assign T663 = wb_reg_sret ? 2'h3 : T664;
  assign T664 = replay_wb ? 2'h2 : 2'h1;

  always @(posedge clk) begin
    wb_reg_xcpt <= T1;
    if(ctrl_killm) begin
      wb_reg_sret <= 1'h0;
    end else begin
      wb_reg_sret <= T5;
    end
    mem_reg_replay <= T7;
    if(ctrl_killx) begin
      mem_reg_replay_next <= 1'h0;
    end else begin
      mem_reg_replay_next <= ex_reg_replay_next;
    end
    if(ctrl_killd) begin
      ex_reg_replay_next <= 1'h0;
    end else begin
      ex_reg_replay_next <= T10;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T79;
    end
    if(ctrl_killd) begin
      ex_reg_mem_val <= 1'h0;
    end else begin
      ex_reg_mem_val <= T88;
    end
    if(reset) begin
      R105 <= 32'h0;
    end else if(T126) begin
      R105 <= T108;
    end else if(io_dpath_ll_wen) begin
      R105 <= T101;
    end
    if(ctrl_killm) begin
      wb_reg_rocc_val <= 1'h0;
    end else begin
      wb_reg_rocc_val <= mem_reg_rocc_val;
    end
    if(ctrl_killx) begin
      mem_reg_rocc_val <= 1'h0;
    end else begin
      mem_reg_rocc_val <= ex_reg_rocc_val;
    end
    if(ctrl_killd) begin
      ex_reg_rocc_val <= 1'h0;
    end else begin
      ex_reg_rocc_val <= T115;
    end
    if(ctrl_killm) begin
      wb_reg_mem_val <= 1'h0;
    end else begin
      wb_reg_mem_val <= mem_reg_mem_val;
    end
    if(ctrl_killx) begin
      mem_reg_mem_val <= 1'h0;
    end else begin
      mem_reg_mem_val <= ex_reg_mem_val;
    end
    if(ctrl_killm) begin
      wb_reg_div_mul_val <= 1'h0;
    end else begin
      wb_reg_div_mul_val <= mem_reg_div_mul_val;
    end
    mem_reg_div_mul_val <= T121;
    if(ctrl_killd) begin
      ex_reg_div_mul_val <= 1'h0;
    end else begin
      ex_reg_div_mul_val <= T123;
    end
    if(ctrl_killm) begin
      wb_reg_fp_val <= 1'h0;
    end else begin
      wb_reg_fp_val <= mem_reg_fp_val;
    end
    if(ctrl_killx) begin
      mem_reg_fp_val <= 1'h0;
    end else begin
      mem_reg_fp_val <= ex_reg_fp_val;
    end
    if(ctrl_killd) begin
      ex_reg_fp_val <= 1'h0;
    end else begin
      ex_reg_fp_val <= 1'h0;
    end
    if(ctrl_killm) begin
      wb_reg_fp_wen <= 1'h0;
    end else begin
      wb_reg_fp_wen <= mem_reg_fp_wen;
    end
    if(ctrl_killx) begin
      mem_reg_fp_wen <= 1'h0;
    end else begin
      mem_reg_fp_wen <= ex_reg_fp_wen;
    end
    if(ctrl_killd) begin
      ex_reg_fp_wen <= 1'h0;
    end else begin
      ex_reg_fp_wen <= 1'h0;
    end
    if(ctrl_killm) begin
      wb_reg_wen <= 1'h0;
    end else begin
      wb_reg_wen <= mem_reg_wen;
    end
    if(ctrl_killx) begin
      mem_reg_wen <= 1'h0;
    end else begin
      mem_reg_wen <= ex_reg_wen;
    end
    if(ctrl_killd) begin
      ex_reg_wen <= 1'h0;
    end else begin
      ex_reg_wen <= id_wen;
    end
    if(T278) begin
      mem_mem_cmd_bh <= ex_slow_bypass;
    end
    if(T246) begin
      ex_reg_mem_type <= T238;
    end
    if(T246) begin
      ex_reg_mem_cmd <= id_mem_cmd;
    end
    if(ctrl_killx) begin
      mem_reg_csr <= 2'h0;
    end else begin
      mem_reg_csr <= ex_reg_csr;
    end
    if(ctrl_killd) begin
      ex_reg_csr <= 2'h0;
    end else begin
      ex_reg_csr <= id_csr;
    end
    if(ctrl_killd) begin
      ex_reg_jalr <= 1'h0;
    end else begin
      ex_reg_jalr <= id_jalr;
    end
    if(ctrl_killx) begin
      mem_reg_jal <= 1'h0;
    end else begin
      mem_reg_jal <= ex_reg_jal;
    end
    if(ctrl_killd) begin
      ex_reg_jal <= 1'h0;
    end else begin
      ex_reg_jal <= id_jal;
    end
    if(ctrl_killx) begin
      mem_reg_jalr <= 1'h0;
    end else begin
      mem_reg_jalr <= ex_reg_jalr;
    end
    if(ctrl_killx) begin
      mem_reg_branch <= 1'h0;
    end else begin
      mem_reg_branch <= ex_reg_branch;
    end
    if(ctrl_killd) begin
      ex_reg_branch <= 1'h0;
    end else begin
      ex_reg_branch <= id_branch;
    end
    if(ctrl_killd) begin
      ex_reg_load_use <= 1'h0;
    end else begin
      ex_reg_load_use <= id_load_use;
    end
    if(ctrl_killx) begin
      mem_reg_sret <= 1'h0;
    end else begin
      mem_reg_sret <= ex_reg_sret;
    end
    if(ctrl_killd) begin
      ex_reg_sret <= 1'h0;
    end else begin
      ex_reg_sret <= id_sret;
    end
    if(ctrl_killx) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= ex_reg_valid;
    end
    if(ctrl_killd) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= 1'h1;
    end
    if(ctrl_killx) begin
      mem_reg_xcpt <= 1'h0;
    end else begin
      mem_reg_xcpt <= ex_xcpt;
    end
    if(ctrl_killd) begin
      ex_reg_xcpt <= 1'h0;
    end else begin
      ex_reg_xcpt <= id_xcpt;
    end
    ex_reg_xcpt_interrupt <= T449;
    wb_reg_replay <= T457;
    mem_reg_xcpt_interrupt <= T468;
    if(ctrl_killm) begin
      wb_reg_flush_inst <= 1'h0;
    end else begin
      wb_reg_flush_inst <= mem_reg_flush_inst;
    end
    if(ctrl_killx) begin
      mem_reg_flush_inst <= 1'h0;
    end else begin
      mem_reg_flush_inst <= ex_reg_flush_inst;
    end
    if(ctrl_killd) begin
      ex_reg_flush_inst <= 1'h0;
    end else begin
      ex_reg_flush_inst <= id_fence_i;
    end
    if(T486) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T485) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(ctrl_killd) begin
      ex_reg_btb_hit <= 1'h0;
    end else begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T486) begin
      mem_reg_btb_resp_bht_index <= ex_reg_btb_resp_bht_index;
    end
    if(T485) begin
      ex_reg_btb_resp_bht_index <= io_imem_btb_resp_bits_bht_index;
    end
    if(T486) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T485) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T486) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T485) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T486) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T485) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T278) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(ctrl_killm) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= mem_reg_valid;
    end
    if(ctrl_killm) begin
      wb_reg_csr <= 2'h0;
    end else begin
      wb_reg_csr <= mem_reg_csr;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out
);

  wire[63:0] sum;
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[31:0] T5;
  wire[63:0] out64;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T133;
  wire cmp;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[63:0] T25;
  wire T26;
  wire[63:0] T27;
  wire T28;
  wire[63:0] T29;
  wire T30;
  wire[63:0] shout_l;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[62:0] T33;
  wire[63:0] T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire[61:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[59:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  wire[63:0] T44;
  wire[55:0] T45;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[47:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[31:0] T53;
  wire[63:0] T54;
  wire[63:0] T134;
  wire[31:0] T55;
  wire[63:0] T56;
  wire[63:0] T135;
  wire[47:0] T57;
  wire[63:0] T58;
  wire[63:0] T136;
  wire[55:0] T59;
  wire[63:0] T60;
  wire[63:0] T137;
  wire[59:0] T61;
  wire[63:0] T62;
  wire[63:0] T138;
  wire[61:0] T63;
  wire[63:0] T64;
  wire[63:0] T139;
  wire[62:0] T65;
  wire T66;
  wire[63:0] shout_r;
  wire[64:0] T67;
  wire[5:0] shamt;
  wire[5:0] T68;
  wire[4:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire[64:0] T73;
  wire[64:0] T74;
  wire[63:0] shin;
  wire[63:0] T75;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[62:0] T78;
  wire[63:0] T79;
  wire[63:0] T80;
  wire[63:0] T81;
  wire[61:0] T82;
  wire[63:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[59:0] T86;
  wire[63:0] T87;
  wire[63:0] T88;
  wire[63:0] T89;
  wire[55:0] T90;
  wire[63:0] T91;
  wire[63:0] T92;
  wire[63:0] T93;
  wire[47:0] T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire[63:0] T97;
  wire[31:0] T98;
  wire[63:0] T99;
  wire[63:0] T140;
  wire[31:0] T100;
  wire[63:0] T101;
  wire[63:0] T141;
  wire[47:0] T102;
  wire[63:0] T103;
  wire[63:0] T142;
  wire[55:0] T104;
  wire[63:0] T105;
  wire[63:0] T143;
  wire[59:0] T106;
  wire[63:0] T107;
  wire[63:0] T144;
  wire[61:0] T108;
  wire[63:0] T109;
  wire[63:0] T145;
  wire[62:0] T110;
  wire[63:0] shin_r;
  wire[31:0] T111;
  wire[31:0] shin_hi;
  wire[31:0] shin_hi_32;
  wire[31:0] T112;
  wire[31:0] T146;
  wire T113;
  wire T114;
  wire[31:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire[31:0] out_hi;
  wire[31:0] T129;
  wire[31:0] T147;
  wire T130;
  wire[31:0] T131;
  wire T132;


  assign io_adder_out = sum;
  assign sum = io_in1 + T0;
  assign T0 = T2 ? T1 : io_in2;
  assign T1 = 64'h0 - io_in2;
  assign T2 = io_fn[2'h3:2'h3];
  assign io_out = T3;
  assign T3 = T4;
  assign T4 = {out_hi, T5};
  assign T5 = out64[5'h1f:1'h0];
  assign out64 = T126 ? sum : T6;
  assign T6 = T123 ? shout_r : T7;
  assign T7 = T66 ? shout_l : T8;
  assign T8 = T30 ? T29 : T9;
  assign T9 = T28 ? T27 : T10;
  assign T10 = T26 ? T25 : T133;
  assign T133 = {63'h0, cmp};
  assign cmp = T24 ^ T11;
  assign T11 = T22 ? T21 : T12;
  assign T12 = T18 ? T17 : T13;
  assign T13 = T16 ? T15 : T14;
  assign T14 = io_in1[6'h3f:6'h3f];
  assign T15 = io_in2[6'h3f:6'h3f];
  assign T16 = io_fn[1'h1:1'h1];
  assign T17 = sum[6'h3f:6'h3f];
  assign T18 = T20 == T19;
  assign T19 = io_in2[6'h3f:6'h3f];
  assign T20 = io_in1[6'h3f:6'h3f];
  assign T21 = sum == 64'h0;
  assign T22 = T23 ^ 1'h1;
  assign T23 = io_fn[2'h2:2'h2];
  assign T24 = io_fn[1'h0:1'h0];
  assign T25 = io_in1 ^ io_in2;
  assign T26 = io_fn == 4'h4;
  assign T27 = io_in1 | io_in2;
  assign T28 = io_fn == 4'h6;
  assign T29 = io_in1 & io_in2;
  assign T30 = io_fn == 4'h7;
  assign shout_l = T64 | T31;
  assign T31 = T32 & 64'haaaaaaaaaaaaaaaa;
  assign T32 = T33 << 1'h1;
  assign T33 = T34[6'h3e:1'h0];
  assign T34 = T62 | T35;
  assign T35 = T36 & 64'hcccccccccccccccc;
  assign T36 = T37 << 2'h2;
  assign T37 = T38[6'h3d:1'h0];
  assign T38 = T60 | T39;
  assign T39 = T40 & 64'hf0f0f0f0f0f0f0f0;
  assign T40 = T41 << 3'h4;
  assign T41 = T42[6'h3b:1'h0];
  assign T42 = T58 | T43;
  assign T43 = T44 & 64'hff00ff00ff00ff00;
  assign T44 = T45 << 4'h8;
  assign T45 = T46[6'h37:1'h0];
  assign T46 = T56 | T47;
  assign T47 = T48 & 64'hffff0000ffff0000;
  assign T48 = T49 << 5'h10;
  assign T49 = T50[6'h2f:1'h0];
  assign T50 = T54 | T51;
  assign T51 = T52 & 64'hffffffff00000000;
  assign T52 = T53 << 6'h20;
  assign T53 = shout_r[5'h1f:1'h0];
  assign T54 = T134 & 64'hffffffff;
  assign T134 = {32'h0, T55};
  assign T55 = shout_r >> 6'h20;
  assign T56 = T135 & 64'hffff0000ffff;
  assign T135 = {16'h0, T57};
  assign T57 = T50 >> 5'h10;
  assign T58 = T136 & 64'hff00ff00ff00ff;
  assign T136 = {8'h0, T59};
  assign T59 = T46 >> 4'h8;
  assign T60 = T137 & 64'hf0f0f0f0f0f0f0f;
  assign T137 = {4'h0, T61};
  assign T61 = T42 >> 3'h4;
  assign T62 = T138 & 64'h3333333333333333;
  assign T138 = {2'h0, T63};
  assign T63 = T38 >> 2'h2;
  assign T64 = T139 & 64'h5555555555555555;
  assign T139 = {1'h0, T65};
  assign T65 = T34 >> 1'h1;
  assign T66 = io_fn == 4'h1;
  assign shout_r = T67[6'h3f:1'h0];
  assign T67 = $signed(T73) >>> shamt;
  assign shamt = T68;
  assign T68 = {T70, T69};
  assign T69 = io_in2[3'h4:1'h0];
  assign T70 = T72 & T71;
  assign T71 = io_dw == 1'h1;
  assign T72 = io_in2[3'h5:3'h5];
  assign T73 = T74;
  assign T74 = {T120, shin};
  assign shin = T117 ? shin_r : T75;
  assign T75 = T109 | T76;
  assign T76 = T77 & 64'haaaaaaaaaaaaaaaa;
  assign T77 = T78 << 1'h1;
  assign T78 = T79[6'h3e:1'h0];
  assign T79 = T107 | T80;
  assign T80 = T81 & 64'hcccccccccccccccc;
  assign T81 = T82 << 2'h2;
  assign T82 = T83[6'h3d:1'h0];
  assign T83 = T105 | T84;
  assign T84 = T85 & 64'hf0f0f0f0f0f0f0f0;
  assign T85 = T86 << 3'h4;
  assign T86 = T87[6'h3b:1'h0];
  assign T87 = T103 | T88;
  assign T88 = T89 & 64'hff00ff00ff00ff00;
  assign T89 = T90 << 4'h8;
  assign T90 = T91[6'h37:1'h0];
  assign T91 = T101 | T92;
  assign T92 = T93 & 64'hffff0000ffff0000;
  assign T93 = T94 << 5'h10;
  assign T94 = T95[6'h2f:1'h0];
  assign T95 = T99 | T96;
  assign T96 = T97 & 64'hffffffff00000000;
  assign T97 = T98 << 6'h20;
  assign T98 = shin_r[5'h1f:1'h0];
  assign T99 = T140 & 64'hffffffff;
  assign T140 = {32'h0, T100};
  assign T100 = shin_r >> 6'h20;
  assign T101 = T141 & 64'hffff0000ffff;
  assign T141 = {16'h0, T102};
  assign T102 = T95 >> 5'h10;
  assign T103 = T142 & 64'hff00ff00ff00ff;
  assign T142 = {8'h0, T104};
  assign T104 = T91 >> 4'h8;
  assign T105 = T143 & 64'hf0f0f0f0f0f0f0f;
  assign T143 = {4'h0, T106};
  assign T106 = T87 >> 3'h4;
  assign T107 = T144 & 64'h3333333333333333;
  assign T144 = {2'h0, T108};
  assign T108 = T83 >> 2'h2;
  assign T109 = T145 & 64'h5555555555555555;
  assign T145 = {1'h0, T110};
  assign T110 = T79 >> 1'h1;
  assign shin_r = {shin_hi, T111};
  assign T111 = io_in1[5'h1f:1'h0];
  assign shin_hi = T116 ? T115 : shin_hi_32;
  assign shin_hi_32 = T114 ? T112 : 32'h0;
  assign T112 = 32'h0 - T146;
  assign T146 = {31'h0, T113};
  assign T113 = io_in1[5'h1f:5'h1f];
  assign T114 = io_fn[2'h3:2'h3];
  assign T115 = io_in1[6'h3f:6'h20];
  assign T116 = io_dw == 1'h1;
  assign T117 = T119 | T118;
  assign T118 = io_fn == 4'hb;
  assign T119 = io_fn == 4'h5;
  assign T120 = T122 & T121;
  assign T121 = shin[6'h3f:6'h3f];
  assign T122 = io_fn[2'h3:2'h3];
  assign T123 = T125 | T124;
  assign T124 = io_fn == 4'hb;
  assign T125 = io_fn == 4'h5;
  assign T126 = T128 | T127;
  assign T127 = io_fn == 4'ha;
  assign T128 = io_fn == 4'h0;
  assign out_hi = T132 ? T131 : T129;
  assign T129 = 32'h0 - T147;
  assign T147 = {31'h0, T130};
  assign T130 = out64[5'h1f:5'h1f];
  assign T131 = out64[6'h3f:6'h20];
  assign T132 = io_dw == 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T140;
  wire[63:0] negated_remainder;
  wire[63:0] T88;
  wire T10;
  wire T11;
  reg  isMul;
  wire T12;
  wire cmdMul;
  wire T13;
  wire[3:0] T14;
  wire T15;
  wire[3:0] T16;
  wire T17;
  wire T18;
  reg [2:0] state;
  wire[2:0] T141;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  reg  neg_out;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  isHi;
  wire T32;
  wire cmdHi;
  wire T33;
  wire T34;
  wire[3:0] T35;
  wire T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire less;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T40;
  wire[64:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire[64:0] T45;
  wire[63:0] rhs_in;
  wire[31:0] T46;
  wire[31:0] T47;
  wire[31:0] T48;
  wire[31:0] T142;
  wire[31:0] T49;
  wire T50;
  wire rhs_sign;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire rhsSigned;
  wire T55;
  wire[3:0] T56;
  wire[64:0] T57;
  wire T58;
  reg [6:0] count;
  wire[6:0] T59;
  wire[6:0] T60;
  wire[6:0] T61;
  wire[6:0] T62;
  wire[6:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire lhs_sign;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire lhsSigned;
  wire T71;
  wire[3:0] T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire[2:0] T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire[2:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire[129:0] T143;
  wire T89;
  wire[129:0] T144;
  wire[63:0] T90;
  wire T91;
  wire[129:0] T92;
  wire[129:0] T93;
  wire[64:0] T94;
  wire[63:0] T95;
  wire[128:0] T96;
  wire[63:0] T97;
  wire[128:0] T98;
  wire[128:0] T99;
  wire[62:0] T100;
  wire[63:0] T101;
  wire[128:0] T102;
  wire[63:0] T103;
  wire[64:0] T104;
  wire[65:0] T105;
  wire[65:0] T145;
  wire[64:0] T106;
  wire[64:0] T107;
  wire T146;
  wire[65:0] T108;
  wire[1:0] T109;
  wire[1:0] T110;
  wire T111;
  wire[64:0] T112;
  wire[64:0] T113;
  wire[64:0] T114;
  wire T115;
  wire T116;
  wire[129:0] T147;
  wire[128:0] T117;
  wire[64:0] T118;
  wire T119;
  wire[63:0] T120;
  wire[63:0] T121;
  wire[63:0] T122;
  wire[63:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[129:0] T148;
  wire[63:0] lhs_in;
  wire[31:0] T127;
  wire[31:0] T128;
  wire[31:0] T129;
  wire[31:0] T149;
  wire[31:0] T130;
  wire T131;
  wire[63:0] T132;
  wire[31:0] T133;
  wire[31:0] T134;
  wire[31:0] T150;
  wire T135;
  wire T136;
  reg  req_dw;
  wire T137;
  wire T138;
  wire T139;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T136 ? T132 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T148 : T5;
  assign T5 = T124 ? T147 : T6;
  assign T6 = T115 ? T92 : T7;
  assign T7 = T91 ? T144 : T8;
  assign T8 = T89 ? T143 : T9;
  assign T9 = T10 ? T140 : remainder;
  assign T140 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T88;
  assign T88 = remainder[6'h3f:1'h0];
  assign T10 = T18 & T11;
  assign T11 = T17 | isMul;
  assign T12 = T1 ? cmdMul : isMul;
  assign cmdMul = T15 | T13;
  assign T13 = T14 == 4'h8;
  assign T14 = io_req_bits_fn & 4'h8;
  assign T15 = T16 == 4'h0;
  assign T16 = io_req_bits_fn & 4'h4;
  assign T17 = remainder[6'h3f:6'h3f];
  assign T18 = state == 3'h1;
  assign T141 = reset ? 3'h0 : T19;
  assign T19 = T1 ? T84 : T20;
  assign T20 = T82 ? 3'h0 : T21;
  assign T21 = T80 ? T78 : T22;
  assign T22 = T76 ? T75 : T23;
  assign T23 = T91 ? T26 : T24;
  assign T24 = T89 ? 3'h5 : T25;
  assign T25 = T18 ? 3'h2 : state;
  assign T26 = neg_out ? 3'h4 : 3'h5;
  assign T27 = T1 ? T64 : T28;
  assign T28 = T29 ? 1'h0 : neg_out;
  assign T29 = T124 & T30;
  assign T30 = T38 & T31;
  assign T31 = isHi ^ 1'h1;
  assign T32 = T1 ? cmdHi : isHi;
  assign cmdHi = T33 | T13;
  assign T33 = T36 | T34;
  assign T34 = T35 == 4'h2;
  assign T35 = io_req_bits_fn & 4'h2;
  assign T36 = T37 == 4'h1;
  assign T37 = io_req_bits_fn & 4'h5;
  assign T38 = T58 & T39;
  assign T39 = less ^ 1'h1;
  assign less = subtractor[7'h40:7'h40];
  assign subtractor = T57 - divisor;
  assign T40 = T1 ? T45 : T41;
  assign T41 = T42 ? subtractor : divisor;
  assign T42 = T18 & T43;
  assign T43 = T44 | isMul;
  assign T44 = divisor[6'h3f:6'h3f];
  assign T45 = {rhs_sign, rhs_in};
  assign rhs_in = {T47, T46};
  assign T46 = io_req_bits_in2[5'h1f:1'h0];
  assign T47 = T50 ? T49 : T48;
  assign T48 = 32'h0 - T142;
  assign T142 = {31'h0, rhs_sign};
  assign T49 = io_req_bits_in2[6'h3f:6'h20];
  assign T50 = io_req_bits_dw == 1'h1;
  assign rhs_sign = rhsSigned & T51;
  assign T51 = T54 ? T53 : T52;
  assign T52 = io_req_bits_in2[5'h1f:5'h1f];
  assign T53 = io_req_bits_in2[6'h3f:6'h3f];
  assign T54 = io_req_bits_dw == 1'h1;
  assign rhsSigned = T55 | T15;
  assign T55 = T56 == 4'h0;
  assign T56 = io_req_bits_fn & 4'h9;
  assign T57 = remainder[8'h80:7'h40];
  assign T58 = count == 7'h0;
  assign T59 = T1 ? 7'h0 : T60;
  assign T60 = T124 ? T63 : T61;
  assign T61 = T115 ? T62 : count;
  assign T62 = count + 7'h1;
  assign T63 = count + 7'h1;
  assign T64 = T74 & T65;
  assign T65 = cmdHi ? lhs_sign : T66;
  assign T66 = lhs_sign != rhs_sign;
  assign lhs_sign = lhsSigned & T67;
  assign T67 = T70 ? T69 : T68;
  assign T68 = io_req_bits_in1[5'h1f:5'h1f];
  assign T69 = io_req_bits_in1[6'h3f:6'h3f];
  assign T70 = io_req_bits_dw == 1'h1;
  assign lhsSigned = T73 | T71;
  assign T71 = T72 == 4'h0;
  assign T72 = io_req_bits_fn & 4'h3;
  assign T73 = T55 | T15;
  assign T74 = cmdMul ^ 1'h1;
  assign T75 = isHi ? 3'h3 : 3'h5;
  assign T76 = T115 & T77;
  assign T77 = count == 7'h3f;
  assign T78 = isHi ? 3'h3 : T79;
  assign T79 = neg_out ? 3'h4 : 3'h5;
  assign T80 = T124 & T81;
  assign T81 = count == 7'h40;
  assign T82 = T83 | io_kill;
  assign T83 = io_resp_ready & io_resp_valid;
  assign T84 = T85 ? 3'h1 : 3'h2;
  assign T85 = lhs_sign | T86;
  assign T86 = rhs_sign & T87;
  assign T87 = cmdMul ^ 1'h1;
  assign T143 = {66'h0, negated_remainder};
  assign T89 = state == 3'h4;
  assign T144 = {66'h0, T90};
  assign T90 = remainder[8'h80:7'h41];
  assign T91 = state == 3'h3;
  assign T92 = T93;
  assign T93 = {T114, T94};
  assign T94 = {1'h0, T95};
  assign T95 = T96[6'h3f:1'h0];
  assign T96 = {T113, T97};
  assign T97 = T98[6'h3f:1'h0];
  assign T98 = T99;
  assign T99 = {T105, T100};
  assign T100 = T101[6'h3f:1'h1];
  assign T101 = T102[6'h3f:1'h0];
  assign T102 = {T104, T103};
  assign T103 = remainder[6'h3f:1'h0];
  assign T104 = remainder[8'h81:7'h41];
  assign T105 = T108 + T145;
  assign T145 = {T146, T106};
  assign T106 = T107;
  assign T107 = T102[8'h80:7'h40];
  assign T146 = T106[7'h40:7'h40];
  assign T108 = $signed(T112) * $signed(T109);
  assign T109 = T110;
  assign T110 = {1'h0, T111};
  assign T111 = T101[1'h0:1'h0];
  assign T112 = divisor;
  assign T113 = T98[8'h80:7'h40];
  assign T114 = T96 >> 7'h40;
  assign T115 = T116 & isMul;
  assign T116 = state == 3'h2;
  assign T147 = {1'h0, T117};
  assign T117 = {T121, T118};
  assign T118 = {T120, T119};
  assign T119 = less ^ 1'h1;
  assign T120 = remainder[6'h3f:1'h0];
  assign T121 = less ? T123 : T122;
  assign T122 = subtractor[6'h3f:1'h0];
  assign T123 = remainder[7'h7f:7'h40];
  assign T124 = T126 & T125;
  assign T125 = isMul ^ 1'h1;
  assign T126 = state == 3'h2;
  assign T148 = {66'h0, lhs_in};
  assign lhs_in = {T128, T127};
  assign T127 = io_req_bits_in1[5'h1f:1'h0];
  assign T128 = T131 ? T130 : T129;
  assign T129 = 32'h0 - T149;
  assign T149 = {31'h0, lhs_sign};
  assign T130 = io_req_bits_in1[6'h3f:6'h20];
  assign T131 = io_req_bits_dw == 1'h1;
  assign T132 = {T134, T133};
  assign T133 = remainder[5'h1f:1'h0];
  assign T134 = 32'h0 - T150;
  assign T150 = {31'h0, T135};
  assign T135 = remainder[5'h1f:5'h1f];
  assign T136 = req_dw == 1'h0;
  assign T137 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T138;
  assign T138 = state == 3'h5;
  assign io_req_ready = T139;
  assign T139 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T148;
    end else if(T124) begin
      remainder <= T147;
    end else if(T115) begin
      remainder <= T92;
    end else if(T91) begin
      remainder <= T144;
    end else if(T89) begin
      remainder <= T143;
    end else if(T10) begin
      remainder <= T140;
    end
    if(T1) begin
      isMul <= cmdMul;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T84;
    end else if(T82) begin
      state <= 3'h0;
    end else if(T80) begin
      state <= T78;
    end else if(T76) begin
      state <= T75;
    end else if(T91) begin
      state <= T26;
    end else if(T89) begin
      state <= 3'h5;
    end else if(T18) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T64;
    end else if(T29) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= cmdHi;
    end
    if(T1) begin
      divisor <= T45;
    end else if(T42) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T124) begin
      count <= T63;
    end else if(T115) begin
      count <= T62;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [11:0] io_rw_addr,
    input [1:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    output[7:0] io_status_ip,
    output[7:0] io_status_im,
    output[6:0] io_status_zero,
    output io_status_er,
    output io_status_vm,
    output io_status_s64,
    output io_status_u64,
    output io_status_ef,
    output io_status_pei,
    output io_status_ei,
    output io_status_ps,
    output io_status_s,
    output[31:0] io_ptbr,
    output[43:0] io_evec,
    input  io_exception,
    input  io_retire,
    input  io_uarch_counters_15,
    input  io_uarch_counters_14,
    input  io_uarch_counters_13,
    input  io_uarch_counters_12,
    input  io_uarch_counters_11,
    input  io_uarch_counters_10,
    input  io_uarch_counters_9,
    input  io_uarch_counters_8,
    input  io_uarch_counters_7,
    input  io_uarch_counters_6,
    input  io_uarch_counters_5,
    input  io_uarch_counters_4,
    input  io_uarch_counters_3,
    input  io_uarch_counters_2,
    input  io_uarch_counters_1,
    input  io_uarch_counters_0,
    input [63:0] io_cause,
    input  io_badvaddr_wen,
    input [43:0] io_pc,
    input  io_sret,
    output io_fatc,
    output io_replay,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  reg [2:0] reg_frm;
  wire[2:0] T468;
  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T469;
  wire[63:0] wdata;
  reg [63:0] host_pcr_bits_data;
  wire[63:0] T2;
  wire[63:0] T3;
  wire T4;
  wire host_pcr_req_fire;
  wire T5;
  reg  host_pcr_req_valid;
  wire T6;
  wire T7;
  wire cpu_req_valid;
  wire T8;
  wire T9;
  reg [41:0] T10;
  wire[11:0] addr;
  wire[11:0] T470;
  wire[10:0] T12;
  wire[10:0] T471;
  reg [4:0] host_pcr_bits_addr;
  wire[4:0] T13;
  wire wen;
  wire T14;
  reg  host_pcr_bits_rw;
  wire T15;
  wire[63:0] T472;
  wire[58:0] T16;
  wire T17;
  wire T18;
  wire[63:0] T19;
  reg [5:0] R20;
  wire[5:0] T473;
  wire[5:0] T21;
  wire[5:0] T22;
  wire[6:0] T23;
  wire[6:0] T474;
  wire[5:0] T24;
  wire[63:0] T25;
  wire T26;
  wire T27;
  reg [57:0] R28;
  wire[57:0] T475;
  wire[57:0] T29;
  wire[57:0] T30;
  wire[57:0] T31;
  wire T32;
  wire[57:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[43:0] T38;
  wire[43:0] T39;
  reg [43:0] reg_epc;
  wire[43:0] T40;
  wire[43:0] T41;
  wire[43:0] T42;
  wire[43:0] T43;
  wire[43:0] T44;
  wire T45;
  wire T46;
  wire[43:0] T476;
  wire[42:0] T47;
  reg [42:0] reg_evec;
  wire[42:0] T48;
  wire[42:0] T49;
  wire[42:0] T50;
  wire T51;
  wire T52;
  wire T477;
  reg [31:0] reg_ptbr;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T55;
  wire[18:0] T56;
  wire T57;
  wire T58;
  reg  reg_status_s;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  reg  reg_status_ps;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  reg  reg_status_ei;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  reg  reg_status_pei;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg  reg_status_ef;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  reg  reg_status_u64;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg  reg_status_s64;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  reg  reg_status_vm;
  wire T91;
  wire T92;
  wire T93;
  reg  reg_status_er;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  reg [6:0] reg_status_zero;
  wire[6:0] T98;
  wire[6:0] T99;
  wire[6:0] T100;
  wire[6:0] T101;
  reg [7:0] reg_status_im;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[7:0] T104;
  wire[7:0] T105;
  wire[3:0] T106;
  wire[1:0] T107;
  reg  r_irq_ipi;
  wire T478;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire[1:0] T113;
  wire T114;
  reg [63:0] reg_fromhost;
  wire[63:0] T479;
  wire[63:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  reg  r_irq_timer;
  wire T480;
  wire T122;
  wire T123;
  wire T124;
  reg [31:0] reg_compare;
  wire[31:0] T125;
  wire[31:0] T126;
  wire[31:0] T127;
  wire[31:0] T128;
  wire T129;
  wire T130;
  wire[63:0] T131;
  wire[63:0] T132;
  wire[63:0] T133;
  reg [5:0] R134;
  wire[5:0] T481;
  wire[5:0] T135;
  wire[5:0] T136;
  wire[6:0] T137;
  wire[6:0] T482;
  wire T138;
  reg [57:0] R139;
  wire[57:0] T483;
  wire[57:0] T140;
  wire[57:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[63:0] T145;
  wire[63:0] T146;
  wire[63:0] T147;
  reg [5:0] R148;
  wire[5:0] T484;
  wire[5:0] T149;
  wire[5:0] T150;
  wire[6:0] T151;
  wire[6:0] T485;
  wire T152;
  reg [57:0] R153;
  wire[57:0] T486;
  wire[57:0] T154;
  wire[57:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[63:0] T159;
  wire[63:0] T160;
  wire[63:0] T161;
  reg [5:0] R162;
  wire[5:0] T487;
  wire[5:0] T163;
  wire[5:0] T164;
  wire[6:0] T165;
  wire[6:0] T488;
  wire T166;
  reg [57:0] R167;
  wire[57:0] T489;
  wire[57:0] T168;
  wire[57:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire[63:0] T173;
  wire[63:0] T174;
  wire[63:0] T175;
  reg [5:0] R176;
  wire[5:0] T490;
  wire[5:0] T177;
  wire[5:0] T178;
  wire[6:0] T179;
  wire[6:0] T491;
  wire T180;
  reg [57:0] R181;
  wire[57:0] T492;
  wire[57:0] T182;
  wire[57:0] T183;
  wire T184;
  wire T185;
  wire T186;
  wire[63:0] T187;
  wire[63:0] T188;
  wire[63:0] T189;
  reg [5:0] R190;
  wire[5:0] T493;
  wire[5:0] T191;
  wire[5:0] T192;
  wire[6:0] T193;
  wire[6:0] T494;
  wire T194;
  reg [57:0] R195;
  wire[57:0] T495;
  wire[57:0] T196;
  wire[57:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire[63:0] T201;
  wire[63:0] T202;
  wire[63:0] T203;
  reg [5:0] R204;
  wire[5:0] T496;
  wire[5:0] T205;
  wire[5:0] T206;
  wire[6:0] T207;
  wire[6:0] T497;
  wire T208;
  reg [57:0] R209;
  wire[57:0] T498;
  wire[57:0] T210;
  wire[57:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire[63:0] T215;
  wire[63:0] T216;
  wire[63:0] T217;
  reg [5:0] R218;
  wire[5:0] T499;
  wire[5:0] T219;
  wire[5:0] T220;
  wire[6:0] T221;
  wire[6:0] T500;
  wire T222;
  reg [57:0] R223;
  wire[57:0] T501;
  wire[57:0] T224;
  wire[57:0] T225;
  wire T226;
  wire T227;
  wire T228;
  wire[63:0] T229;
  wire[63:0] T230;
  wire[63:0] T231;
  reg [5:0] R232;
  wire[5:0] T502;
  wire[5:0] T233;
  wire[5:0] T234;
  wire[6:0] T235;
  wire[6:0] T503;
  wire T236;
  reg [57:0] R237;
  wire[57:0] T504;
  wire[57:0] T238;
  wire[57:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[63:0] T243;
  wire[63:0] T244;
  wire[63:0] T245;
  reg [5:0] R246;
  wire[5:0] T505;
  wire[5:0] T247;
  wire[5:0] T248;
  wire[6:0] T249;
  wire[6:0] T506;
  wire T250;
  reg [57:0] R251;
  wire[57:0] T507;
  wire[57:0] T252;
  wire[57:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire[63:0] T257;
  wire[63:0] T258;
  wire[63:0] T259;
  reg [5:0] R260;
  wire[5:0] T508;
  wire[5:0] T261;
  wire[5:0] T262;
  wire[6:0] T263;
  wire[6:0] T509;
  wire T264;
  reg [57:0] R265;
  wire[57:0] T510;
  wire[57:0] T266;
  wire[57:0] T267;
  wire T268;
  wire T269;
  wire T270;
  wire[63:0] T271;
  wire[63:0] T272;
  wire[63:0] T273;
  reg [5:0] R274;
  wire[5:0] T511;
  wire[5:0] T275;
  wire[5:0] T276;
  wire[6:0] T277;
  wire[6:0] T512;
  wire T278;
  reg [57:0] R279;
  wire[57:0] T513;
  wire[57:0] T280;
  wire[57:0] T281;
  wire T282;
  wire T283;
  wire T284;
  wire[63:0] T285;
  wire[63:0] T286;
  wire[63:0] T287;
  reg [5:0] R288;
  wire[5:0] T514;
  wire[5:0] T289;
  wire[5:0] T290;
  wire[6:0] T291;
  wire[6:0] T515;
  wire T292;
  reg [57:0] R293;
  wire[57:0] T516;
  wire[57:0] T294;
  wire[57:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[63:0] T299;
  wire[63:0] T300;
  wire[63:0] T301;
  reg [5:0] R302;
  wire[5:0] T517;
  wire[5:0] T303;
  wire[5:0] T304;
  wire[6:0] T305;
  wire[6:0] T518;
  wire T306;
  reg [57:0] R307;
  wire[57:0] T519;
  wire[57:0] T308;
  wire[57:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[63:0] T313;
  wire[63:0] T314;
  wire[63:0] T315;
  reg [5:0] R316;
  wire[5:0] T520;
  wire[5:0] T317;
  wire[5:0] T318;
  wire[6:0] T319;
  wire[6:0] T521;
  wire T320;
  reg [57:0] R321;
  wire[57:0] T522;
  wire[57:0] T322;
  wire[57:0] T323;
  wire T324;
  wire T325;
  wire T326;
  wire[63:0] T327;
  wire[63:0] T328;
  wire[63:0] T329;
  reg [5:0] R330;
  wire[5:0] T523;
  wire[5:0] T331;
  wire[5:0] T332;
  wire[6:0] T333;
  wire[6:0] T524;
  wire T334;
  reg [57:0] R335;
  wire[57:0] T525;
  wire[57:0] T336;
  wire[57:0] T337;
  wire T338;
  wire T339;
  wire T340;
  wire[63:0] T341;
  wire[63:0] T342;
  wire[63:0] T343;
  reg [5:0] R344;
  wire[5:0] T526;
  wire[5:0] T345;
  wire[5:0] T346;
  wire[6:0] T347;
  wire[6:0] T527;
  wire T348;
  reg [57:0] R349;
  wire[57:0] T528;
  wire[57:0] T350;
  wire[57:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[63:0] T355;
  wire[63:0] T356;
  wire[63:0] T357;
  wire[63:0] T358;
  reg [63:0] reg_tohost;
  wire[63:0] T529;
  wire[63:0] T359;
  wire[63:0] T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire[63:0] T369;
  wire[63:0] T530;
  wire T370;
  reg  reg_stats;
  wire T531;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire[63:0] T375;
  wire[63:0] T532;
  wire[1:0] T376;
  wire[63:0] T377;
  wire[63:0] T533;
  wire[1:0] T378;
  wire T379;
  wire[63:0] T380;
  wire[63:0] T534;
  wire[1:0] T381;
  wire[63:0] T382;
  wire[63:0] T535;
  wire[1:0] T383;
  wire T384;
  wire[63:0] T385;
  wire[63:0] T536;
  wire T386;
  wire T387;
  wire[63:0] T388;
  wire[63:0] T537;
  wire[31:0] T389;
  wire[31:0] T390;
  wire[31:0] T391;
  wire[5:0] T392;
  wire[2:0] T393;
  wire[1:0] T394;
  wire[2:0] T395;
  wire[1:0] T396;
  wire[25:0] T397;
  wire[2:0] T398;
  wire[1:0] T399;
  wire[22:0] T400;
  wire[14:0] T401;
  wire[63:0] T402;
  wire[63:0] T403;
  reg [63:0] reg_cause;
  wire[63:0] T404;
  wire T405;
  wire[63:0] T406;
  wire[63:0] T538;
  wire[42:0] T407;
  wire[63:0] T408;
  wire[63:0] T539;
  wire[31:0] T409;
  wire[63:0] T410;
  wire[63:0] T411;
  wire[63:0] T412;
  wire[63:0] T413;
  wire[63:0] T540;
  wire[31:0] T414;
  wire[31:0] read_ptbr;
  wire[18:0] T415;
  wire[63:0] T416;
  wire[63:0] T541;
  wire[42:0] T417;
  reg [42:0] reg_badvaddr;
  wire[42:0] T542;
  wire[43:0] T418;
  wire[43:0] T543;
  wire[43:0] T419;
  wire[43:0] T420;
  wire[42:0] T421;
  wire T422;
  wire T423;
  wire[20:0] T424;
  wire T425;
  wire T426;
  wire[42:0] T427;
  wire T428;
  wire[63:0] T429;
  wire[63:0] T544;
  wire[43:0] T430;
  wire[63:0] T431;
  wire[63:0] T432;
  reg [63:0] reg_sup1;
  wire[63:0] T433;
  wire T434;
  wire T435;
  wire[63:0] T436;
  wire[63:0] T437;
  reg [63:0] reg_sup0;
  wire[63:0] T438;
  wire T439;
  wire T440;
  wire[63:0] T441;
  wire[63:0] T442;
  wire[63:0] T443;
  reg [5:0] R444;
  wire[5:0] T545;
  wire[5:0] T445;
  wire[5:0] T446;
  wire[6:0] T447;
  wire[6:0] T546;
  wire T448;
  reg [57:0] R449;
  wire[57:0] T547;
  wire[57:0] T450;
  wire[57:0] T451;
  wire T452;
  wire T453;
  wire T454;
  wire[63:0] T455;
  wire[63:0] T456;
  wire T457;
  wire[63:0] T458;
  wire[63:0] T459;
  wire T460;
  wire T548;
  wire T461;
  reg  host_pcr_rep_valid;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    reg_frm = {1{$random}};
    host_pcr_bits_data = {2{$random}};
    host_pcr_req_valid = {1{$random}};
    host_pcr_bits_addr = {1{$random}};
    host_pcr_bits_rw = {1{$random}};
    R20 = {1{$random}};
    R28 = {2{$random}};
    reg_epc = {2{$random}};
    reg_evec = {2{$random}};
    reg_ptbr = {1{$random}};
    reg_status_s = {1{$random}};
    reg_status_ps = {1{$random}};
    reg_status_ei = {1{$random}};
    reg_status_pei = {1{$random}};
    reg_status_ef = {1{$random}};
    reg_status_u64 = {1{$random}};
    reg_status_s64 = {1{$random}};
    reg_status_vm = {1{$random}};
    reg_status_er = {1{$random}};
    reg_status_zero = {1{$random}};
    reg_status_im = {1{$random}};
    r_irq_ipi = {1{$random}};
    reg_fromhost = {2{$random}};
    r_irq_timer = {1{$random}};
    reg_compare = {1{$random}};
    R134 = {1{$random}};
    R139 = {2{$random}};
    R148 = {1{$random}};
    R153 = {2{$random}};
    R162 = {1{$random}};
    R167 = {2{$random}};
    R176 = {1{$random}};
    R181 = {2{$random}};
    R190 = {1{$random}};
    R195 = {2{$random}};
    R204 = {1{$random}};
    R209 = {2{$random}};
    R218 = {1{$random}};
    R223 = {2{$random}};
    R232 = {1{$random}};
    R237 = {2{$random}};
    R246 = {1{$random}};
    R251 = {2{$random}};
    R260 = {1{$random}};
    R265 = {2{$random}};
    R274 = {1{$random}};
    R279 = {2{$random}};
    R288 = {1{$random}};
    R293 = {2{$random}};
    R302 = {1{$random}};
    R307 = {2{$random}};
    R316 = {1{$random}};
    R321 = {2{$random}};
    R330 = {1{$random}};
    R335 = {2{$random}};
    R344 = {1{$random}};
    R349 = {2{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_cause = {2{$random}};
    reg_badvaddr = {2{$random}};
    reg_sup1 = {2{$random}};
    reg_sup0 = {2{$random}};
    R444 = {1{$random}};
    R449 = {2{$random}};
    host_pcr_rep_valid = {1{$random}};
  end
`endif

  assign io_fcsr_rm = reg_frm;
  assign T468 = T0[2'h2:1'h0];
  assign T0 = T17 ? T472 : T1;
  assign T1 = T8 ? wdata : T469;
  assign T469 = {61'h0, reg_frm};
  assign wdata = cpu_req_valid ? io_rw_wdata : host_pcr_bits_data;
  assign T2 = host_pcr_req_fire ? io_rw_rdata : T3;
  assign T3 = T4 ? io_host_pcr_req_bits_data : host_pcr_bits_data;
  assign T4 = io_host_pcr_req_ready & io_host_pcr_req_valid;
  assign host_pcr_req_fire = host_pcr_req_valid & T5;
  assign T5 = cpu_req_valid ^ 1'h1;
  assign T6 = host_pcr_req_fire ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : host_pcr_req_valid;
  assign cpu_req_valid = io_rw_cmd != 2'h0;
  assign T8 = wen & T9;
  assign T9 = T10[1'h1:1'h1];
  always @(*) case (addr)
    1: T10 = 42'h1;
    2: T10 = 42'h2;
    3: T10 = 42'h4;
    192: T10 = 42'h8;
    1280: T10 = 42'h10;
    1281: T10 = 42'h20;
    1282: T10 = 42'h40;
    1283: T10 = 42'h80;
    1284: T10 = 42'h100;
    1285: T10 = 42'h200;
    1286: T10 = 42'h400;
    1287: T10 = 42'h800;
    1288: T10 = 42'h1000;
    1289: T10 = 42'h2000;
    1290: T10 = 42'h4000;
    1291: T10 = 42'h8000;
    1292: T10 = 42'h10000;
    1293: T10 = 42'h20000;
    1294: T10 = 42'h40000;
    1295: T10 = 42'h80000;
    1309: T10 = 42'h100000;
    1310: T10 = 42'h200000;
    1311: T10 = 42'h400000;
    3072: T10 = 42'h800000;
    3073: T10 = 42'h1000000;
    3074: T10 = 42'h2000000;
    3264: T10 = 42'h4000000;
    3265: T10 = 42'h8000000;
    3266: T10 = 42'h10000000;
    3267: T10 = 42'h20000000;
    3268: T10 = 42'h40000000;
    3269: T10 = 42'h80000000;
    3270: T10 = 42'h100000000;
    3271: T10 = 42'h200000000;
    3272: T10 = 42'h400000000;
    3273: T10 = 42'h800000000;
    3274: T10 = 42'h1000000000;
    3275: T10 = 42'h2000000000;
    3276: T10 = 42'h4000000000;
    3277: T10 = 42'h8000000000;
    3278: T10 = 42'h10000000000;
    3279: T10 = 42'h20000000000;
`ifndef SYNTHESIS
    default: T10 = {2{$random}};
`else
    default: T10 = 42'bx;
`endif
  endcase
  assign addr = cpu_req_valid ? io_rw_addr : T470;
  assign T470 = {1'h0, T12};
  assign T12 = T471 | 11'h500;
  assign T471 = {6'h0, host_pcr_bits_addr};
  assign T13 = T4 ? io_host_pcr_req_bits_addr : host_pcr_bits_addr;
  assign wen = cpu_req_valid | T14;
  assign T14 = host_pcr_req_fire & host_pcr_bits_rw;
  assign T15 = T4 ? io_host_pcr_req_bits_rw : host_pcr_bits_rw;
  assign T472 = {5'h0, T16};
  assign T16 = wdata >> 3'h5;
  assign T17 = wen & T18;
  assign T18 = T10[2'h2:2'h2];
  assign io_time = T19;
  assign T19 = {R28, R20};
  assign T473 = reset ? 6'h0 : T21;
  assign T21 = T26 ? T24 : T22;
  assign T22 = T23[3'h5:1'h0];
  assign T23 = T474 + 7'h1;
  assign T474 = {1'h0, R20};
  assign T24 = T25[3'h5:1'h0];
  assign T25 = wdata;
  assign T26 = wen & T27;
  assign T27 = T10[4'ha:4'ha];
  assign T475 = reset ? 58'h0 : T29;
  assign T29 = T26 ? T33 : T30;
  assign T30 = T32 ? T31 : R28;
  assign T31 = R28 + 58'h1;
  assign T32 = T23[3'h6:3'h6];
  assign T33 = T25[6'h3f:3'h6];
  assign io_replay = T34;
  assign T34 = io_host_ipi_req_valid & T35;
  assign T35 = io_host_ipi_req_ready ^ 1'h1;
  assign io_fatc = T36;
  assign T36 = wen & T37;
  assign T37 = T10[5'h11:5'h11];
  assign io_evec = T38;
  assign T38 = T39;
  assign T39 = io_exception ? T476 : reg_epc;
  assign T40 = T45 ? T43 : T41;
  assign T41 = io_exception ? T42 : reg_epc;
  assign T42 = io_pc;
  assign T43 = T44;
  assign T44 = wdata[6'h2b:1'h0];
  assign T45 = wen & T46;
  assign T46 = T10[3'h6:3'h6];
  assign T476 = {T477, T47};
  assign T47 = reg_evec;
  assign T48 = T51 ? T49 : reg_evec;
  assign T49 = T50;
  assign T50 = wdata[6'h2a:1'h0];
  assign T51 = wen & T52;
  assign T52 = T10[4'hc:4'hc];
  assign T477 = T47[6'h2a:6'h2a];
  assign io_ptbr = reg_ptbr;
  assign T53 = T57 ? T54 : reg_ptbr;
  assign T54 = T55;
  assign T55 = {T56, 13'h0};
  assign T56 = wdata[5'h1f:4'hd];
  assign T57 = wen & T58;
  assign T58 = T10[4'h8:4'h8];
  assign io_status_s = reg_status_s;
  assign T59 = reset ? 1'h1 : T60;
  assign T60 = T68 ? T67 : T61;
  assign T61 = io_sret ? reg_status_ps : T62;
  assign T62 = io_exception ? 1'h1 : reg_status_s;
  assign T63 = reset ? 1'h0 : T64;
  assign T64 = T68 ? T66 : T65;
  assign T65 = io_exception ? reg_status_s : reg_status_ps;
  assign T66 = wdata[1'h1:1'h1];
  assign T67 = wdata[1'h0:1'h0];
  assign T68 = wen & T69;
  assign T69 = T10[4'he:4'he];
  assign io_status_ps = reg_status_ps;
  assign io_status_ei = reg_status_ei;
  assign T70 = reset ? 1'h0 : T71;
  assign T71 = T68 ? T78 : T72;
  assign T72 = io_sret ? reg_status_pei : T73;
  assign T73 = io_exception ? 1'h0 : reg_status_ei;
  assign T74 = reset ? 1'h0 : T75;
  assign T75 = T68 ? T77 : T76;
  assign T76 = io_exception ? reg_status_ei : reg_status_pei;
  assign T77 = wdata[2'h3:2'h3];
  assign T78 = wdata[2'h2:2'h2];
  assign io_status_pei = reg_status_pei;
  assign io_status_ef = reg_status_ef;
  assign T79 = reset ? 1'h0 : T80;
  assign T80 = T68 ? 1'h0 : T81;
  assign T81 = T68 ? T82 : reg_status_ef;
  assign T82 = wdata[3'h4:3'h4];
  assign io_status_u64 = reg_status_u64;
  assign T83 = reset ? 1'h1 : T84;
  assign T84 = T68 ? 1'h1 : T85;
  assign T85 = T68 ? T86 : reg_status_u64;
  assign T86 = wdata[3'h5:3'h5];
  assign io_status_s64 = reg_status_s64;
  assign T87 = reset ? 1'h1 : T88;
  assign T88 = T68 ? 1'h1 : T89;
  assign T89 = T68 ? T90 : reg_status_s64;
  assign T90 = wdata[3'h6:3'h6];
  assign io_status_vm = reg_status_vm;
  assign T91 = reset ? 1'h0 : T92;
  assign T92 = T68 ? T93 : reg_status_vm;
  assign T93 = wdata[3'h7:3'h7];
  assign io_status_er = reg_status_er;
  assign T94 = reset ? 1'h0 : T95;
  assign T95 = T68 ? 1'h0 : T96;
  assign T96 = T68 ? T97 : reg_status_er;
  assign T97 = wdata[4'h8:4'h8];
  assign io_status_zero = reg_status_zero;
  assign T98 = reset ? 7'h0 : T99;
  assign T99 = T68 ? 7'h0 : T100;
  assign T100 = T68 ? T101 : reg_status_zero;
  assign T101 = wdata[4'hf:4'h9];
  assign io_status_im = reg_status_im;
  assign T102 = reset ? 8'h0 : T103;
  assign T103 = T68 ? T104 : reg_status_im;
  assign T104 = wdata[5'h17:5'h10];
  assign io_status_ip = T105;
  assign T105 = {T106, 4'h0};
  assign T106 = {T113, T107};
  assign T107 = {r_irq_ipi, 1'h0};
  assign T478 = reset ? 1'h1 : T108;
  assign T108 = io_host_ipi_rep_valid ? 1'h1 : T109;
  assign T109 = T111 ? T110 : r_irq_ipi;
  assign T110 = wdata[1'h0:1'h0];
  assign T111 = wen & T112;
  assign T112 = T10[5'h13:5'h13];
  assign T113 = {r_irq_timer, T114};
  assign T114 = reg_fromhost != 64'h0;
  assign T479 = reset ? 64'h0 : T115;
  assign T115 = T116 ? wdata : reg_fromhost;
  assign T116 = T120 & T117;
  assign T117 = T119 | T118;
  assign T118 = host_pcr_req_fire ^ 1'h1;
  assign T119 = reg_fromhost == 64'h0;
  assign T120 = wen & T121;
  assign T121 = T10[5'h16:5'h16];
  assign T480 = reset ? 1'h0 : T122;
  assign T122 = T129 ? 1'h0 : T123;
  assign T123 = T124 ? 1'h1 : r_irq_timer;
  assign T124 = T128 == reg_compare;
  assign T125 = T129 ? T126 : reg_compare;
  assign T126 = T127;
  assign T127 = wdata[5'h1f:1'h0];
  assign T128 = T19[5'h1f:1'h0];
  assign T129 = wen & T130;
  assign T130 = T10[4'hb:4'hb];
  assign io_rw_rdata = T131;
  assign T131 = T145 | T132;
  assign T132 = T144 ? T133 : 64'h0;
  assign T133 = {R139, R134};
  assign T481 = reset ? 6'h0 : T135;
  assign T135 = T138 ? T136 : R134;
  assign T136 = T137[3'h5:1'h0];
  assign T137 = T482 + 7'h1;
  assign T482 = {1'h0, R134};
  assign T138 = io_uarch_counters_15 != 1'h0;
  assign T483 = reset ? 58'h0 : T140;
  assign T140 = T142 ? T141 : R139;
  assign T141 = R139 + 58'h1;
  assign T142 = T138 & T143;
  assign T143 = T137[3'h6:3'h6];
  assign T144 = T10[6'h29:6'h29];
  assign T145 = T159 | T146;
  assign T146 = T158 ? T147 : 64'h0;
  assign T147 = {R153, R148};
  assign T484 = reset ? 6'h0 : T149;
  assign T149 = T152 ? T150 : R148;
  assign T150 = T151[3'h5:1'h0];
  assign T151 = T485 + 7'h1;
  assign T485 = {1'h0, R148};
  assign T152 = io_uarch_counters_14 != 1'h0;
  assign T486 = reset ? 58'h0 : T154;
  assign T154 = T156 ? T155 : R153;
  assign T155 = R153 + 58'h1;
  assign T156 = T152 & T157;
  assign T157 = T151[3'h6:3'h6];
  assign T158 = T10[6'h28:6'h28];
  assign T159 = T173 | T160;
  assign T160 = T172 ? T161 : 64'h0;
  assign T161 = {R167, R162};
  assign T487 = reset ? 6'h0 : T163;
  assign T163 = T166 ? T164 : R162;
  assign T164 = T165[3'h5:1'h0];
  assign T165 = T488 + 7'h1;
  assign T488 = {1'h0, R162};
  assign T166 = io_uarch_counters_13 != 1'h0;
  assign T489 = reset ? 58'h0 : T168;
  assign T168 = T170 ? T169 : R167;
  assign T169 = R167 + 58'h1;
  assign T170 = T166 & T171;
  assign T171 = T165[3'h6:3'h6];
  assign T172 = T10[6'h27:6'h27];
  assign T173 = T187 | T174;
  assign T174 = T186 ? T175 : 64'h0;
  assign T175 = {R181, R176};
  assign T490 = reset ? 6'h0 : T177;
  assign T177 = T180 ? T178 : R176;
  assign T178 = T179[3'h5:1'h0];
  assign T179 = T491 + 7'h1;
  assign T491 = {1'h0, R176};
  assign T180 = io_uarch_counters_12 != 1'h0;
  assign T492 = reset ? 58'h0 : T182;
  assign T182 = T184 ? T183 : R181;
  assign T183 = R181 + 58'h1;
  assign T184 = T180 & T185;
  assign T185 = T179[3'h6:3'h6];
  assign T186 = T10[6'h26:6'h26];
  assign T187 = T201 | T188;
  assign T188 = T200 ? T189 : 64'h0;
  assign T189 = {R195, R190};
  assign T493 = reset ? 6'h0 : T191;
  assign T191 = T194 ? T192 : R190;
  assign T192 = T193[3'h5:1'h0];
  assign T193 = T494 + 7'h1;
  assign T494 = {1'h0, R190};
  assign T194 = io_uarch_counters_11 != 1'h0;
  assign T495 = reset ? 58'h0 : T196;
  assign T196 = T198 ? T197 : R195;
  assign T197 = R195 + 58'h1;
  assign T198 = T194 & T199;
  assign T199 = T193[3'h6:3'h6];
  assign T200 = T10[6'h25:6'h25];
  assign T201 = T215 | T202;
  assign T202 = T214 ? T203 : 64'h0;
  assign T203 = {R209, R204};
  assign T496 = reset ? 6'h0 : T205;
  assign T205 = T208 ? T206 : R204;
  assign T206 = T207[3'h5:1'h0];
  assign T207 = T497 + 7'h1;
  assign T497 = {1'h0, R204};
  assign T208 = io_uarch_counters_10 != 1'h0;
  assign T498 = reset ? 58'h0 : T210;
  assign T210 = T212 ? T211 : R209;
  assign T211 = R209 + 58'h1;
  assign T212 = T208 & T213;
  assign T213 = T207[3'h6:3'h6];
  assign T214 = T10[6'h24:6'h24];
  assign T215 = T229 | T216;
  assign T216 = T228 ? T217 : 64'h0;
  assign T217 = {R223, R218};
  assign T499 = reset ? 6'h0 : T219;
  assign T219 = T222 ? T220 : R218;
  assign T220 = T221[3'h5:1'h0];
  assign T221 = T500 + 7'h1;
  assign T500 = {1'h0, R218};
  assign T222 = io_uarch_counters_9 != 1'h0;
  assign T501 = reset ? 58'h0 : T224;
  assign T224 = T226 ? T225 : R223;
  assign T225 = R223 + 58'h1;
  assign T226 = T222 & T227;
  assign T227 = T221[3'h6:3'h6];
  assign T228 = T10[6'h23:6'h23];
  assign T229 = T243 | T230;
  assign T230 = T242 ? T231 : 64'h0;
  assign T231 = {R237, R232};
  assign T502 = reset ? 6'h0 : T233;
  assign T233 = T236 ? T234 : R232;
  assign T234 = T235[3'h5:1'h0];
  assign T235 = T503 + 7'h1;
  assign T503 = {1'h0, R232};
  assign T236 = io_uarch_counters_8 != 1'h0;
  assign T504 = reset ? 58'h0 : T238;
  assign T238 = T240 ? T239 : R237;
  assign T239 = R237 + 58'h1;
  assign T240 = T236 & T241;
  assign T241 = T235[3'h6:3'h6];
  assign T242 = T10[6'h22:6'h22];
  assign T243 = T257 | T244;
  assign T244 = T256 ? T245 : 64'h0;
  assign T245 = {R251, R246};
  assign T505 = reset ? 6'h0 : T247;
  assign T247 = T250 ? T248 : R246;
  assign T248 = T249[3'h5:1'h0];
  assign T249 = T506 + 7'h1;
  assign T506 = {1'h0, R246};
  assign T250 = io_uarch_counters_7 != 1'h0;
  assign T507 = reset ? 58'h0 : T252;
  assign T252 = T254 ? T253 : R251;
  assign T253 = R251 + 58'h1;
  assign T254 = T250 & T255;
  assign T255 = T249[3'h6:3'h6];
  assign T256 = T10[6'h21:6'h21];
  assign T257 = T271 | T258;
  assign T258 = T270 ? T259 : 64'h0;
  assign T259 = {R265, R260};
  assign T508 = reset ? 6'h0 : T261;
  assign T261 = T264 ? T262 : R260;
  assign T262 = T263[3'h5:1'h0];
  assign T263 = T509 + 7'h1;
  assign T509 = {1'h0, R260};
  assign T264 = io_uarch_counters_6 != 1'h0;
  assign T510 = reset ? 58'h0 : T266;
  assign T266 = T268 ? T267 : R265;
  assign T267 = R265 + 58'h1;
  assign T268 = T264 & T269;
  assign T269 = T263[3'h6:3'h6];
  assign T270 = T10[6'h20:6'h20];
  assign T271 = T285 | T272;
  assign T272 = T284 ? T273 : 64'h0;
  assign T273 = {R279, R274};
  assign T511 = reset ? 6'h0 : T275;
  assign T275 = T278 ? T276 : R274;
  assign T276 = T277[3'h5:1'h0];
  assign T277 = T512 + 7'h1;
  assign T512 = {1'h0, R274};
  assign T278 = io_uarch_counters_5 != 1'h0;
  assign T513 = reset ? 58'h0 : T280;
  assign T280 = T282 ? T281 : R279;
  assign T281 = R279 + 58'h1;
  assign T282 = T278 & T283;
  assign T283 = T277[3'h6:3'h6];
  assign T284 = T10[5'h1f:5'h1f];
  assign T285 = T299 | T286;
  assign T286 = T298 ? T287 : 64'h0;
  assign T287 = {R293, R288};
  assign T514 = reset ? 6'h0 : T289;
  assign T289 = T292 ? T290 : R288;
  assign T290 = T291[3'h5:1'h0];
  assign T291 = T515 + 7'h1;
  assign T515 = {1'h0, R288};
  assign T292 = io_uarch_counters_4 != 1'h0;
  assign T516 = reset ? 58'h0 : T294;
  assign T294 = T296 ? T295 : R293;
  assign T295 = R293 + 58'h1;
  assign T296 = T292 & T297;
  assign T297 = T291[3'h6:3'h6];
  assign T298 = T10[5'h1e:5'h1e];
  assign T299 = T313 | T300;
  assign T300 = T312 ? T301 : 64'h0;
  assign T301 = {R307, R302};
  assign T517 = reset ? 6'h0 : T303;
  assign T303 = T306 ? T304 : R302;
  assign T304 = T305[3'h5:1'h0];
  assign T305 = T518 + 7'h1;
  assign T518 = {1'h0, R302};
  assign T306 = io_uarch_counters_3 != 1'h0;
  assign T519 = reset ? 58'h0 : T308;
  assign T308 = T310 ? T309 : R307;
  assign T309 = R307 + 58'h1;
  assign T310 = T306 & T311;
  assign T311 = T305[3'h6:3'h6];
  assign T312 = T10[5'h1d:5'h1d];
  assign T313 = T327 | T314;
  assign T314 = T326 ? T315 : 64'h0;
  assign T315 = {R321, R316};
  assign T520 = reset ? 6'h0 : T317;
  assign T317 = T320 ? T318 : R316;
  assign T318 = T319[3'h5:1'h0];
  assign T319 = T521 + 7'h1;
  assign T521 = {1'h0, R316};
  assign T320 = io_uarch_counters_2 != 1'h0;
  assign T522 = reset ? 58'h0 : T322;
  assign T322 = T324 ? T323 : R321;
  assign T323 = R321 + 58'h1;
  assign T324 = T320 & T325;
  assign T325 = T319[3'h6:3'h6];
  assign T326 = T10[5'h1c:5'h1c];
  assign T327 = T341 | T328;
  assign T328 = T340 ? T329 : 64'h0;
  assign T329 = {R335, R330};
  assign T523 = reset ? 6'h0 : T331;
  assign T331 = T334 ? T332 : R330;
  assign T332 = T333[3'h5:1'h0];
  assign T333 = T524 + 7'h1;
  assign T524 = {1'h0, R330};
  assign T334 = io_uarch_counters_1 != 1'h0;
  assign T525 = reset ? 58'h0 : T336;
  assign T336 = T338 ? T337 : R335;
  assign T337 = R335 + 58'h1;
  assign T338 = T334 & T339;
  assign T339 = T333[3'h6:3'h6];
  assign T340 = T10[5'h1b:5'h1b];
  assign T341 = T355 | T342;
  assign T342 = T354 ? T343 : 64'h0;
  assign T343 = {R349, R344};
  assign T526 = reset ? 6'h0 : T345;
  assign T345 = T348 ? T346 : R344;
  assign T346 = T347[3'h5:1'h0];
  assign T347 = T527 + 7'h1;
  assign T527 = {1'h0, R344};
  assign T348 = io_uarch_counters_0 != 1'h0;
  assign T528 = reset ? 58'h0 : T350;
  assign T350 = T352 ? T351 : R349;
  assign T351 = R349 + 58'h1;
  assign T352 = T348 & T353;
  assign T353 = T347[3'h6:3'h6];
  assign T354 = T10[5'h1a:5'h1a];
  assign T355 = T357 | T356;
  assign T356 = T121 ? reg_fromhost : 64'h0;
  assign T357 = T369 | T358;
  assign T358 = T368 ? reg_tohost : 64'h0;
  assign T529 = reset ? 64'h0 : T359;
  assign T359 = T364 ? wdata : T360;
  assign T360 = T361 ? 64'h0 : reg_tohost;
  assign T361 = T362 & T368;
  assign T362 = host_pcr_req_fire & T363;
  assign T363 = host_pcr_bits_rw ^ 1'h1;
  assign T364 = T367 & T365;
  assign T365 = T366 | host_pcr_req_fire;
  assign T366 = reg_tohost == 64'h0;
  assign T367 = wen & T368;
  assign T368 = T10[5'h15:5'h15];
  assign T369 = T375 | T530;
  assign T530 = {63'h0, T370};
  assign T370 = T374 ? reg_stats : 1'h0;
  assign T531 = reset ? 1'h0 : T371;
  assign T371 = T373 ? T372 : reg_stats;
  assign T372 = wdata[1'h0:1'h0];
  assign T373 = wen & T374;
  assign T374 = T10[2'h3:2'h3];
  assign T375 = T377 | T532;
  assign T532 = {62'h0, T376};
  assign T376 = T112 ? 2'h2 : 2'h0;
  assign T377 = T380 | T533;
  assign T533 = {62'h0, T378};
  assign T378 = T379 ? 2'h2 : 2'h0;
  assign T379 = T10[5'h12:5'h12];
  assign T380 = T382 | T534;
  assign T534 = {62'h0, T381};
  assign T381 = T37 ? 2'h2 : 2'h0;
  assign T382 = T385 | T535;
  assign T535 = {62'h0, T383};
  assign T383 = T384 ? 2'h2 : 2'h0;
  assign T384 = T10[5'h10:5'h10];
  assign T385 = T388 | T536;
  assign T536 = {63'h0, T386};
  assign T386 = T387 ? io_host_id : 1'h0;
  assign T387 = T10[4'hf:4'hf];
  assign T388 = T402 | T537;
  assign T537 = {32'h0, T389};
  assign T389 = T69 ? T390 : 32'h0;
  assign T390 = T391;
  assign T391 = {T397, T392};
  assign T392 = {T395, T393};
  assign T393 = {io_status_ei, T394};
  assign T394 = {io_status_ps, io_status_s};
  assign T395 = {io_status_u64, T396};
  assign T396 = {io_status_ef, io_status_pei};
  assign T397 = {T400, T398};
  assign T398 = {io_status_er, T399};
  assign T399 = {io_status_vm, io_status_s64};
  assign T400 = {io_status_ip, T401};
  assign T401 = {io_status_im, io_status_zero};
  assign T402 = T406 | T403;
  assign T403 = T405 ? reg_cause : 64'h0;
  assign T404 = io_exception ? io_cause : reg_cause;
  assign T405 = T10[4'hd:4'hd];
  assign T406 = T408 | T538;
  assign T538 = {21'h0, T407};
  assign T407 = T52 ? reg_evec : 43'h0;
  assign T408 = T410 | T539;
  assign T539 = {32'h0, T409};
  assign T409 = T130 ? reg_compare : 32'h0;
  assign T410 = T412 | T411;
  assign T411 = T27 ? T19 : 64'h0;
  assign T412 = T413 | 64'h0;
  assign T413 = T416 | T540;
  assign T540 = {32'h0, T414};
  assign T414 = T58 ? read_ptbr : 32'h0;
  assign read_ptbr = T415 << 4'hd;
  assign T415 = reg_ptbr[5'h1f:4'hd];
  assign T416 = T429 | T541;
  assign T541 = {21'h0, T417};
  assign T417 = T428 ? reg_badvaddr : 43'h0;
  assign T542 = T418[6'h2a:1'h0];
  assign T418 = io_badvaddr_wen ? T419 : T543;
  assign T543 = {1'h0, reg_badvaddr};
  assign T419 = T420;
  assign T420 = {T422, T421};
  assign T421 = io_rw_wdata[6'h2a:1'h0];
  assign T422 = T426 ? T425 : T423;
  assign T423 = T424 != 21'h0;
  assign T424 = io_rw_wdata[6'h3f:6'h2b];
  assign T425 = T424 == 21'h1fffff;
  assign T426 = $signed(T427) < $signed(1'h0);
  assign T427 = T421;
  assign T428 = T10[3'h7:3'h7];
  assign T429 = T431 | T544;
  assign T544 = {20'h0, T430};
  assign T430 = T46 ? reg_epc : 44'h0;
  assign T431 = T436 | T432;
  assign T432 = T435 ? reg_sup1 : 64'h0;
  assign T433 = T434 ? wdata : reg_sup1;
  assign T434 = wen & T435;
  assign T435 = T10[3'h5:3'h5];
  assign T436 = T441 | T437;
  assign T437 = T440 ? reg_sup0 : 64'h0;
  assign T438 = T439 ? wdata : reg_sup0;
  assign T439 = wen & T440;
  assign T440 = T10[3'h4:3'h4];
  assign T441 = T455 | T442;
  assign T442 = T454 ? T443 : 64'h0;
  assign T443 = {R449, R444};
  assign T545 = reset ? 6'h0 : T445;
  assign T445 = T448 ? T446 : R444;
  assign T446 = T447[3'h5:1'h0];
  assign T447 = T546 + 7'h1;
  assign T546 = {1'h0, R444};
  assign T448 = io_retire != 1'h0;
  assign T547 = reset ? 58'h0 : T450;
  assign T450 = T452 ? T451 : R449;
  assign T451 = R449 + 58'h1;
  assign T452 = T448 & T453;
  assign T453 = T447[3'h6:3'h6];
  assign T454 = T10[5'h19:5'h19];
  assign T455 = T458 | T456;
  assign T456 = T457 ? T19 : 64'h0;
  assign T457 = T10[5'h18:5'h18];
  assign T458 = 64'h0 | T459;
  assign T459 = T460 ? T19 : 64'h0;
  assign T460 = T10[5'h17:5'h17];
  assign io_host_debug_stats_pcr = reg_stats;
  assign io_host_ipi_rep_ready = 1'h1;
  assign io_host_ipi_req_bits = T548;
  assign T548 = io_rw_wdata[1'h0:1'h0];
  assign io_host_ipi_req_valid = T461;
  assign T461 = cpu_req_valid & T379;
  assign io_host_pcr_rep_bits = host_pcr_bits_data;
  assign io_host_pcr_rep_valid = host_pcr_rep_valid;
  assign T462 = T464 ? 1'h0 : T463;
  assign T463 = host_pcr_req_fire ? 1'h1 : host_pcr_rep_valid;
  assign T464 = io_host_pcr_rep_ready & io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = T465;
  assign T465 = T467 & T466;
  assign T466 = host_pcr_rep_valid ^ 1'h1;
  assign T467 = host_pcr_req_valid ^ 1'h1;

  always @(posedge clk) begin
    reg_frm <= T468;
    if(host_pcr_req_fire) begin
      host_pcr_bits_data <= io_rw_rdata;
    end else if(T4) begin
      host_pcr_bits_data <= io_host_pcr_req_bits_data;
    end
    if(host_pcr_req_fire) begin
      host_pcr_req_valid <= 1'h0;
    end else if(T4) begin
      host_pcr_req_valid <= 1'h1;
    end
    if(T4) begin
      host_pcr_bits_addr <= io_host_pcr_req_bits_addr;
    end
    if(T4) begin
      host_pcr_bits_rw <= io_host_pcr_req_bits_rw;
    end
    if(reset) begin
      R20 <= 6'h0;
    end else if(T26) begin
      R20 <= T24;
    end else begin
      R20 <= T22;
    end
    if(reset) begin
      R28 <= 58'h0;
    end else if(T26) begin
      R28 <= T33;
    end else if(T32) begin
      R28 <= T31;
    end
    if(T45) begin
      reg_epc <= T43;
    end else if(io_exception) begin
      reg_epc <= T42;
    end
    if(T51) begin
      reg_evec <= T49;
    end
    if(T57) begin
      reg_ptbr <= T54;
    end
    if(reset) begin
      reg_status_s <= 1'h1;
    end else if(T68) begin
      reg_status_s <= T67;
    end else if(io_sret) begin
      reg_status_s <= reg_status_ps;
    end else if(io_exception) begin
      reg_status_s <= 1'h1;
    end
    if(reset) begin
      reg_status_ps <= 1'h0;
    end else if(T68) begin
      reg_status_ps <= T66;
    end else if(io_exception) begin
      reg_status_ps <= reg_status_s;
    end
    if(reset) begin
      reg_status_ei <= 1'h0;
    end else if(T68) begin
      reg_status_ei <= T78;
    end else if(io_sret) begin
      reg_status_ei <= reg_status_pei;
    end else if(io_exception) begin
      reg_status_ei <= 1'h0;
    end
    if(reset) begin
      reg_status_pei <= 1'h0;
    end else if(T68) begin
      reg_status_pei <= T77;
    end else if(io_exception) begin
      reg_status_pei <= reg_status_ei;
    end
    if(reset) begin
      reg_status_ef <= 1'h0;
    end else if(T68) begin
      reg_status_ef <= 1'h0;
    end else if(T68) begin
      reg_status_ef <= T82;
    end
    if(reset) begin
      reg_status_u64 <= 1'h1;
    end else if(T68) begin
      reg_status_u64 <= 1'h1;
    end else if(T68) begin
      reg_status_u64 <= T86;
    end
    if(reset) begin
      reg_status_s64 <= 1'h1;
    end else if(T68) begin
      reg_status_s64 <= 1'h1;
    end else if(T68) begin
      reg_status_s64 <= T90;
    end
    if(reset) begin
      reg_status_vm <= 1'h0;
    end else if(T68) begin
      reg_status_vm <= T93;
    end
    if(reset) begin
      reg_status_er <= 1'h0;
    end else if(T68) begin
      reg_status_er <= 1'h0;
    end else if(T68) begin
      reg_status_er <= T97;
    end
    if(reset) begin
      reg_status_zero <= 7'h0;
    end else if(T68) begin
      reg_status_zero <= 7'h0;
    end else if(T68) begin
      reg_status_zero <= T101;
    end
    if(reset) begin
      reg_status_im <= 8'h0;
    end else if(T68) begin
      reg_status_im <= T104;
    end
    if(reset) begin
      r_irq_ipi <= 1'h1;
    end else if(io_host_ipi_rep_valid) begin
      r_irq_ipi <= 1'h1;
    end else if(T111) begin
      r_irq_ipi <= T110;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T116) begin
      reg_fromhost <= wdata;
    end
    if(reset) begin
      r_irq_timer <= 1'h0;
    end else if(T129) begin
      r_irq_timer <= 1'h0;
    end else if(T124) begin
      r_irq_timer <= 1'h1;
    end
    if(T129) begin
      reg_compare <= T126;
    end
    if(reset) begin
      R134 <= 6'h0;
    end else if(T138) begin
      R134 <= T136;
    end
    if(reset) begin
      R139 <= 58'h0;
    end else if(T142) begin
      R139 <= T141;
    end
    if(reset) begin
      R148 <= 6'h0;
    end else if(T152) begin
      R148 <= T150;
    end
    if(reset) begin
      R153 <= 58'h0;
    end else if(T156) begin
      R153 <= T155;
    end
    if(reset) begin
      R162 <= 6'h0;
    end else if(T166) begin
      R162 <= T164;
    end
    if(reset) begin
      R167 <= 58'h0;
    end else if(T170) begin
      R167 <= T169;
    end
    if(reset) begin
      R176 <= 6'h0;
    end else if(T180) begin
      R176 <= T178;
    end
    if(reset) begin
      R181 <= 58'h0;
    end else if(T184) begin
      R181 <= T183;
    end
    if(reset) begin
      R190 <= 6'h0;
    end else if(T194) begin
      R190 <= T192;
    end
    if(reset) begin
      R195 <= 58'h0;
    end else if(T198) begin
      R195 <= T197;
    end
    if(reset) begin
      R204 <= 6'h0;
    end else if(T208) begin
      R204 <= T206;
    end
    if(reset) begin
      R209 <= 58'h0;
    end else if(T212) begin
      R209 <= T211;
    end
    if(reset) begin
      R218 <= 6'h0;
    end else if(T222) begin
      R218 <= T220;
    end
    if(reset) begin
      R223 <= 58'h0;
    end else if(T226) begin
      R223 <= T225;
    end
    if(reset) begin
      R232 <= 6'h0;
    end else if(T236) begin
      R232 <= T234;
    end
    if(reset) begin
      R237 <= 58'h0;
    end else if(T240) begin
      R237 <= T239;
    end
    if(reset) begin
      R246 <= 6'h0;
    end else if(T250) begin
      R246 <= T248;
    end
    if(reset) begin
      R251 <= 58'h0;
    end else if(T254) begin
      R251 <= T253;
    end
    if(reset) begin
      R260 <= 6'h0;
    end else if(T264) begin
      R260 <= T262;
    end
    if(reset) begin
      R265 <= 58'h0;
    end else if(T268) begin
      R265 <= T267;
    end
    if(reset) begin
      R274 <= 6'h0;
    end else if(T278) begin
      R274 <= T276;
    end
    if(reset) begin
      R279 <= 58'h0;
    end else if(T282) begin
      R279 <= T281;
    end
    if(reset) begin
      R288 <= 6'h0;
    end else if(T292) begin
      R288 <= T290;
    end
    if(reset) begin
      R293 <= 58'h0;
    end else if(T296) begin
      R293 <= T295;
    end
    if(reset) begin
      R302 <= 6'h0;
    end else if(T306) begin
      R302 <= T304;
    end
    if(reset) begin
      R307 <= 58'h0;
    end else if(T310) begin
      R307 <= T309;
    end
    if(reset) begin
      R316 <= 6'h0;
    end else if(T320) begin
      R316 <= T318;
    end
    if(reset) begin
      R321 <= 58'h0;
    end else if(T324) begin
      R321 <= T323;
    end
    if(reset) begin
      R330 <= 6'h0;
    end else if(T334) begin
      R330 <= T332;
    end
    if(reset) begin
      R335 <= 58'h0;
    end else if(T338) begin
      R335 <= T337;
    end
    if(reset) begin
      R344 <= 6'h0;
    end else if(T348) begin
      R344 <= T346;
    end
    if(reset) begin
      R349 <= 58'h0;
    end else if(T352) begin
      R349 <= T351;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T364) begin
      reg_tohost <= wdata;
    end else if(T361) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T373) begin
      reg_stats <= T372;
    end
    if(io_exception) begin
      reg_cause <= io_cause;
    end
    reg_badvaddr <= T542;
    if(T434) begin
      reg_sup1 <= wdata;
    end
    if(T439) begin
      reg_sup0 <= wdata;
    end
    if(reset) begin
      R444 <= 6'h0;
    end else if(T448) begin
      R444 <= T446;
    end
    if(reset) begin
      R449 <= 58'h0;
    end else if(T452) begin
      R449 <= T451;
    end
    if(T464) begin
      host_pcr_rep_valid <= 1'h0;
    end else if(host_pcr_req_fire) begin
      host_pcr_rep_valid <= 1'h1;
    end
  end
endmodule

module Datapath(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [2:0] io_ctrl_sel_pc,
    input  io_ctrl_killd,
    input  io_ctrl_ren_1,
    input  io_ctrl_ren_0,
    input [2:0] io_ctrl_sel_alu2,
    input [1:0] io_ctrl_sel_alu1,
    input [2:0] io_ctrl_sel_imm,
    input  io_ctrl_fn_dw,
    input [3:0] io_ctrl_fn_alu,
    input  io_ctrl_div_mul_val,
    input  io_ctrl_div_mul_kill,
    //input  io_ctrl_div_val
    //input  io_ctrl_div_kill
    input [2:0] io_ctrl_csr,
    input  io_ctrl_sret,
    input  io_ctrl_mem_load,
    input  io_ctrl_wb_load,
    input  io_ctrl_ex_fp_val,
    input  io_ctrl_mem_fp_val,
    input  io_ctrl_ex_wen,
    input  io_ctrl_ex_valid,
    input  io_ctrl_mem_jalr,
    input  io_ctrl_mem_branch,
    input  io_ctrl_mem_wen,
    input  io_ctrl_wb_wen,
    input [2:0] io_ctrl_ex_mem_type,
    input  io_ctrl_ex_rs2_val,
    input  io_ctrl_ex_rocc_val,
    input  io_ctrl_mem_rocc_val,
    input  io_ctrl_bypass_1,
    input  io_ctrl_bypass_0,
    input [1:0] io_ctrl_bypass_src_1,
    input [1:0] io_ctrl_bypass_src_0,
    input  io_ctrl_ll_ready,
    input  io_ctrl_retire,
    input  io_ctrl_exception,
    input [63:0] io_ctrl_cause,
    input  io_ctrl_badvaddr_wen,
    output[31:0] io_ctrl_inst,
    //output io_ctrl_jalr_eq
    output io_ctrl_mem_br_taken,
    output io_ctrl_mem_misprediction,
    output io_ctrl_div_mul_rdy,
    output io_ctrl_ll_wen,
    output[4:0] io_ctrl_ll_waddr,
    output[4:0] io_ctrl_ex_waddr,
    output io_ctrl_mem_rs1_ra,
    output[4:0] io_ctrl_mem_waddr,
    output[4:0] io_ctrl_wb_waddr,
    output[7:0] io_ctrl_status_ip,
    output[7:0] io_ctrl_status_im,
    output[6:0] io_ctrl_status_zero,
    output io_ctrl_status_er,
    output io_ctrl_status_vm,
    output io_ctrl_status_s64,
    output io_ctrl_status_u64,
    output io_ctrl_status_ef,
    output io_ctrl_status_pei,
    output io_ctrl_status_ei,
    output io_ctrl_status_ps,
    output io_ctrl_status_s,
    output io_ctrl_fp_sboard_clr,
    output[4:0] io_ctrl_fp_sboard_clra,
    output io_ctrl_csr_replay,
    input  io_dmem_req_ready,
    //output io_dmem_req_valid
    //output io_dmem_req_bits_kill
    //output[2:0] io_dmem_req_bits_typ
    //output io_dmem_req_bits_phys
    output[43:0] io_dmem_req_bits_addr,
    output[63:0] io_dmem_req_bits_data,
    output[7:0] io_dmem_req_bits_tag,
    //output[4:0] io_dmem_req_bits_cmd
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    //output io_imem_req_valid
    output[43:0] io_imem_req_bits_pc,
    //output io_imem_resp_ready
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_index,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    //output io_imem_btb_update_valid
    //output io_imem_btb_update_bits_prediction_valid
    //output io_imem_btb_update_bits_prediction_bits_taken
    //output[42:0] io_imem_btb_update_bits_prediction_bits_target
    //output[2:0] io_imem_btb_update_bits_prediction_bits_entry
    //output[3:0] io_imem_btb_update_bits_prediction_bits_bht_index
    //output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    //output io_imem_btb_update_bits_taken
    //output io_imem_btb_update_bits_isJump
    //output io_imem_btb_update_bits_isCall
    //output io_imem_btb_update_bits_isReturn
    //output io_imem_btb_update_bits_incorrectTarget
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    //output io_imem_invalidate
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  reg  ex_reg_kill;
  wire T7;
  reg  mem_reg_kill;
  wire[31:0] T8;
  wire[63:0] T9;
  reg [63:0] R10;
  reg [63:0] R11;
  wire[63:0] ex_rs_1;
  wire[63:0] T12;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[63:0] id_rs_1;
  wire[63:0] T16;
  wire[63:0] T17;
  reg [63:0] T18 [30:0];
  wire[63:0] T19;
  wire T20;
  wire T21;
  wire[4:0] T22;
  wire T23;
  wire T24;
  wire[4:0] wb_waddr;
  wire wb_wen;
  wire[4:0] T25;
  wire[4:0] T26;
  wire[4:0] T27;
  wire[63:0] wb_wdata;
  wire[63:0] T28;
  wire[63:0] T29;
  wire[63:0] T30;
  reg [63:0] wb_reg_wdata;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[63:0] mem_int_wdata;
  reg [63:0] mem_reg_wdata;
  wire[63:0] T33;
  wire[63:0] T200;
  wire[44:0] mem_br_target;
  wire[44:0] T34;
  wire[44:0] T35;
  reg [43:0] mem_reg_pc;
  wire[43:0] T36;
  reg [43:0] ex_reg_pc;
  wire[43:0] T37;
  wire[44:0] T201;
  wire[21:0] T38;
  wire[21:0] T39;
  wire[21:0] T40;
  wire[21:0] T41;
  wire[11:0] T42;
  wire[4:0] T43;
  wire[3:0] T44;
  wire[6:0] T45;
  wire[5:0] T46;
  wire T47;
  wire T48;
  wire[9:0] T49;
  wire[8:0] T50;
  wire[7:0] T51;
  wire[7:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[21:0] T202;
  wire[14:0] T58;
  wire[14:0] T59;
  wire[11:0] T60;
  wire[4:0] T61;
  wire[3:0] T62;
  wire[6:0] T63;
  wire[5:0] T64;
  wire T65;
  wire T66;
  wire[2:0] T67;
  wire[1:0] T68;
  wire T69;
  wire T70;
  wire[6:0] T203;
  wire T204;
  wire T71;
  wire[22:0] T205;
  wire T206;
  wire[18:0] T207;
  wire T208;
  wire T72;
  wire T73;
  wire[63:0] ll_wdata;
  wire T74;
  wire dmem_resp_xpu;
  wire T75;
  wire T76;
  wire dmem_resp_valid;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T81;
  wire[61:0] T82;
  wire T83;
  wire T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[63:0] T209;
  wire bypass_0;
  wire[63:0] bypass_1;
  wire T87;
  wire[1:0] T88;
  wire[63:0] T89;
  wire[63:0] bypass_2;
  wire[63:0] bypass_3;
  wire T90;
  wire T91;
  reg  ex_reg_rs_bypass_1;
  wire T92;
  wire[4:0] T93;
  wire[4:0] T94;
  wire[63:0] T95;
  reg [63:0] R96;
  reg [63:0] R97;
  wire[63:0] ex_rs_0;
  wire[63:0] T98;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T99;
  wire[1:0] T100;
  wire[1:0] T101;
  wire[63:0] id_rs_0;
  wire[63:0] T102;
  wire[63:0] T103;
  wire[4:0] T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T110;
  wire[61:0] T111;
  wire T112;
  wire T113;
  wire[63:0] T114;
  wire[63:0] T115;
  wire[63:0] T210;
  wire T116;
  wire[1:0] T117;
  wire[63:0] T118;
  wire T119;
  wire T120;
  reg  ex_reg_rs_bypass_0;
  wire T121;
  wire[4:0] T122;
  wire[4:0] T123;
  wire T124;
  wire[63:0] T125;
  wire[4:0] T126;
  wire[4:0] T127;
  wire[43:0] T128;
  reg [43:0] wb_reg_pc;
  wire[43:0] T129;
  wire T130;
  wire[32:0] T131;
  wire[32:0] T132;
  wire T133;
  wire[1135:0] T134;
  wire[63:0] T223;
  wire[63:0] T224;
  wire[63:0] T225;
  wire[63:0] T226;
  wire T227;
  wire[63:0] T228;
  wire T229;
  wire[1:0] T230;
  wire[11:0] T231;
  wire T232;
  wire T193;
  wire dmem_resp_replay;
  reg  ex_reg_ctrl_fn_dw;
  wire T233;
  wire T234;
  reg [3:0] ex_reg_ctrl_fn_alu;
  wire[3:0] T235;
  wire[63:0] ex_op1;
  wire[63:0] T236;
  wire[43:0] T237;
  wire[43:0] T238;
  wire T239;
  reg [1:0] ex_reg_sel_alu1;
  wire[1:0] T240;
  wire[19:0] T241;
  wire T242;
  wire[63:0] T243;
  wire T244;
  wire[63:0] T245;
  wire[63:0] ex_op2;
  wire[63:0] T246;
  wire[31:0] T247;
  wire[31:0] T248;
  wire[3:0] T249;
  wire T250;
  reg [2:0] ex_reg_sel_alu2;
  wire[2:0] T251;
  wire[27:0] T252;
  wire T253;
  wire[31:0] ex_imm;
  wire[31:0] T254;
  wire[11:0] T255;
  wire[4:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  reg [2:0] ex_reg_sel_imm;
  wire[2:0] T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[3:0] T270;
  wire[3:0] T271;
  wire T272;
  wire[3:0] T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire[6:0] T278;
  wire[5:0] T279;
  wire[5:0] T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[19:0] T298;
  wire[18:0] T299;
  wire[7:0] T300;
  wire[7:0] T301;
  wire[7:0] T302;
  wire[7:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[10:0] T307;
  wire[10:0] T308;
  wire[10:0] T309;
  wire[10:0] T310;
  wire T311;
  wire T312;
  wire[31:0] T313;
  wire T314;
  wire[63:0] T315;
  wire T316;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T135;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T136;
  wire[6:0] T137;
  wire[4:0] T138;
  wire T139;
  wire T140;
  wire T141;
  wire[4:0] T142;
  wire[4:0] T143;
  wire[6:0] T144;
  wire[4:0] T211;
  wire[6:0] dmem_resp_waddr;
  wire[7:0] T145;
  wire T146;
  wire dmem_resp_fpu;
  wire T147;
  wire[42:0] T212;
  wire[42:0] T213;
  wire[42:0] T214;
  wire[43:0] T215;
  wire[44:0] T148;
  wire[44:0] T149;
  wire[44:0] T216;
  wire[43:0] T150;
  wire T151;
  wire[44:0] mem_npc;
  wire[44:0] T217;
  wire[43:0] T152;
  wire[42:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire[1:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire[21:0] T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire[7:0] T218;
  wire[5:0] T168;
  wire[63:0] T169;
  wire[43:0] T170;
  wire[43:0] T171;
  wire[42:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire[1:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire[21:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[4:0] T219;
  wire T186;
  wire[4:0] T187;
  wire[4:0] T188;
  wire T189;
  wire[4:0] T190;
  wire[4:0] T191;
  wire[4:0] T220;
  wire[6:0] T192;
  wire[6:0] T221;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire[44:0] T222;
  wire T199;
  wire[63:0] alu_io_out;
  wire[63:0] alu_io_adder_out;
  wire div_io_req_ready;
  wire div_io_resp_valid;
  wire[63:0] div_io_resp_bits_data;
  wire[4:0] div_io_resp_bits_tag;
  wire pcr_io_host_pcr_req_ready;
  wire pcr_io_host_pcr_rep_valid;
  wire[63:0] pcr_io_host_pcr_rep_bits;
  wire pcr_io_host_ipi_req_valid;
  wire pcr_io_host_ipi_req_bits;
  wire pcr_io_host_ipi_rep_ready;
  wire pcr_io_host_debug_stats_pcr;
  wire[63:0] pcr_io_rw_rdata;
  wire[7:0] pcr_io_status_ip;
  wire[7:0] pcr_io_status_im;
  wire[6:0] pcr_io_status_zero;
  wire pcr_io_status_er;
  wire pcr_io_status_vm;
  wire pcr_io_status_s64;
  wire pcr_io_status_u64;
  wire pcr_io_status_ef;
  wire pcr_io_status_pei;
  wire pcr_io_status_ei;
  wire pcr_io_status_ps;
  wire pcr_io_status_s;
  wire[31:0] pcr_io_ptbr;
  wire[43:0] pcr_io_evec;
  wire pcr_io_fatc;
  wire pcr_io_replay;
  wire[63:0] pcr_io_time;
  wire[2:0] pcr_io_fcsr_rm;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    ex_reg_kill = {1{$random}};
    mem_reg_kill = {1{$random}};
    R10 = {2{$random}};
    R11 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T18[initvar] = {2{$random}};
    wb_reg_wdata = {2{$random}};
    mem_reg_wdata = {2{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R96 = {2{$random}};
    R97 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    ex_reg_ctrl_fn_dw = {1{$random}};
    ex_reg_ctrl_fn_alu = {1{$random}};
    ex_reg_sel_alu1 = {1{$random}};
    ex_reg_sel_alu2 = {1{$random}};
    ex_reg_sel_imm = {1{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
  end
`endif

  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T7 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T6 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data : ex_reg_inst;
  assign T5 = io_ctrl_killd ^ 1'h1;
  assign T6 = ex_reg_kill ^ 1'h1;
  assign T7 = mem_reg_kill ^ 1'h1;
  assign T8 = wb_reg_inst;
  assign T9 = R10;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T85 : T12;
  assign T12 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T13 = T80 ? io_ctrl_bypass_src_1 : T14;
  assign T14 = T79 ? T15 : ex_reg_rs_lsb_1;
  assign T15 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T16;
  assign T16 = T77 ? wb_wdata : T17;
  assign T17 = T18[T26];
  assign T20 = T23 & T21;
  assign T21 = T22 < 5'h1f;
  assign T22 = T25[3'h4:1'h0];
  assign T23 = wb_wen & T24;
  assign T24 = wb_waddr != 5'h0;
  assign wb_waddr = io_ctrl_ll_wen ? io_ctrl_ll_waddr : io_ctrl_wb_waddr;
  assign wb_wen = io_ctrl_ll_wen | io_ctrl_wb_wen;
  assign T25 = ~ wb_waddr;
  assign T26 = ~ T27;
  assign T27 = io_imem_resp_bits_data[5'h18:5'h14];
  assign wb_wdata = T28;
  assign T28 = T74 ? io_dmem_resp_bits_data_subword : T29;
  assign T29 = io_ctrl_ll_wen ? ll_wdata : T30;
  assign T30 = T73 ? pcr_io_rw_rdata : wb_reg_wdata;
  assign T31 = T7 ? T32 : wb_reg_wdata;
  assign T32 = T72 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = io_ctrl_mem_jalr ? T200 : mem_reg_wdata;
  assign T33 = T6 ? alu_io_out : mem_reg_wdata;
  assign T200 = {T207, mem_br_target};
  assign mem_br_target = T201 + T34;
  assign T34 = T35;
  assign T35 = {1'h0, mem_reg_pc};
  assign T36 = T6 ? ex_reg_pc : mem_reg_pc;
  assign T37 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T201 = {T205, T38};
  assign T38 = T71 ? T202 : T39;
  assign T39 = T55 ? T40 : 22'h4;
  assign T40 = T41;
  assign T41 = {T49, T42};
  assign T42 = {T45, T43};
  assign T43 = {T44, 1'h0};
  assign T44 = mem_reg_inst[5'h18:5'h15];
  assign T45 = {T47, T46};
  assign T46 = mem_reg_inst[5'h1e:5'h19];
  assign T47 = T48;
  assign T48 = mem_reg_inst[5'h14:5'h14];
  assign T49 = {T53, T50};
  assign T50 = {T53, T51};
  assign T51 = T52;
  assign T52 = mem_reg_inst[5'h13:4'hc];
  assign T53 = T54;
  assign T54 = mem_reg_inst[5'h1f:5'h1f];
  assign T55 = T57 & T56;
  assign T56 = io_ctrl_mem_branch ^ 1'h1;
  assign T57 = io_ctrl_mem_jalr ^ 1'h1;
  assign T202 = {T203, T58};
  assign T58 = T59;
  assign T59 = {T67, T60};
  assign T60 = {T63, T61};
  assign T61 = {T62, 1'h0};
  assign T62 = mem_reg_inst[4'hb:4'h8];
  assign T63 = {T65, T64};
  assign T64 = mem_reg_inst[5'h1e:5'h19];
  assign T65 = T66;
  assign T66 = mem_reg_inst[3'h7:3'h7];
  assign T67 = {T69, T68};
  assign T68 = {T69, T69};
  assign T69 = T70;
  assign T70 = mem_reg_inst[5'h1f:5'h1f];
  assign T203 = T204 ? 7'h7f : 7'h0;
  assign T204 = T58[4'he:4'he];
  assign T71 = io_ctrl_mem_branch & io_ctrl_mem_br_taken;
  assign T205 = T206 ? 23'h7fffff : 23'h0;
  assign T206 = T38[5'h15:5'h15];
  assign T207 = T208 ? 19'h7ffff : 19'h0;
  assign T208 = mem_br_target[6'h2c:6'h2c];
  assign T72 = io_ctrl_mem_fp_val & io_ctrl_mem_wen;
  assign T73 = io_ctrl_csr != 3'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign T74 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_xpu = T75 ^ 1'h1;
  assign T75 = T76;
  assign T76 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T77 = T23 & T78;
  assign T78 = wb_waddr == T27;
  assign T79 = T5 & io_ctrl_ren_1;
  assign T80 = T5 & io_ctrl_bypass_1;
  assign T81 = T83 ? T82 : ex_reg_rs_msb_1;
  assign T82 = id_rs_1 >> 2'h2;
  assign T83 = T79 & T84;
  assign T84 = io_ctrl_bypass_1 ^ 1'h1;
  assign T85 = T91 ? T89 : T86;
  assign T86 = T87 ? bypass_1 : T209;
  assign T209 = {63'h0, bypass_0};
  assign bypass_0 = 1'h0;
  assign bypass_1 = mem_reg_wdata;
  assign T87 = T88[1'h0:1'h0];
  assign T88 = ex_reg_rs_lsb_1;
  assign T89 = T90 ? bypass_3 : bypass_2;
  assign bypass_2 = wb_reg_wdata;
  assign bypass_3 = io_dmem_resp_bits_data;
  assign T90 = T88[1'h0:1'h0];
  assign T91 = T88[1'h1:1'h1];
  assign T92 = T5 ? io_ctrl_bypass_1 : ex_reg_rs_bypass_1;
  assign T93 = T94;
  assign T94 = wb_reg_inst[5'h18:5'h14];
  assign T95 = R96;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T114 : T98;
  assign T98 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T99 = T109 ? io_ctrl_bypass_src_0 : T100;
  assign T100 = T108 ? T101 : ex_reg_rs_lsb_0;
  assign T101 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T102;
  assign T102 = T106 ? wb_wdata : T103;
  assign T103 = T18[T104];
  assign T104 = ~ T105;
  assign T105 = io_imem_resp_bits_data[5'h13:4'hf];
  assign T106 = T23 & T107;
  assign T107 = wb_waddr == T105;
  assign T108 = T5 & io_ctrl_ren_0;
  assign T109 = T5 & io_ctrl_bypass_0;
  assign T110 = T112 ? T111 : ex_reg_rs_msb_0;
  assign T111 = id_rs_0 >> 2'h2;
  assign T112 = T108 & T113;
  assign T113 = io_ctrl_bypass_0 ^ 1'h1;
  assign T114 = T120 ? T118 : T115;
  assign T115 = T116 ? bypass_1 : T210;
  assign T210 = {63'h0, bypass_0};
  assign T116 = T117[1'h0:1'h0];
  assign T117 = ex_reg_rs_lsb_0;
  assign T118 = T119 ? bypass_3 : bypass_2;
  assign T119 = T117[1'h0:1'h0];
  assign T120 = T117[1'h1:1'h1];
  assign T121 = T5 ? io_ctrl_bypass_0 : ex_reg_rs_bypass_0;
  assign T122 = T123;
  assign T123 = wb_reg_inst[5'h13:4'hf];
  assign T124 = wb_wen;
  assign T125 = wb_wdata;
  assign T126 = T127;
  assign T127 = wb_wen ? wb_waddr : 5'h0;
  assign T128 = wb_reg_pc;
  assign T129 = T7 ? mem_reg_pc : wb_reg_pc;
  assign T130 = io_ctrl_retire;
  assign T131 = T132;
  assign T132 = pcr_io_time[6'h20:1'h0];
  assign T133 = io_host_id;
  assign T223 = T229 ? T228 : T224;
  assign T224 = T227 ? T225 : wb_reg_wdata;
  assign T225 = pcr_io_rw_rdata & T226;
  assign T226 = ~ wb_reg_wdata;
  assign T227 = io_ctrl_csr == 3'h3;
  assign T228 = pcr_io_rw_rdata | wb_reg_wdata;
  assign T229 = io_ctrl_csr == 3'h2;
  assign T230 = io_ctrl_csr[1'h1:1'h0];
  assign T231 = wb_reg_inst[5'h1f:5'h14];
  assign T232 = T193 ? 1'h0 : io_ctrl_ll_ready;
  assign T193 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign T233 = T5 ? T234 : ex_reg_ctrl_fn_dw;
  assign T234 = io_ctrl_fn_dw;
  assign T235 = T5 ? io_ctrl_fn_alu : ex_reg_ctrl_fn_alu;
  assign ex_op1 = T244 ? T243 : T236;
  assign T236 = {T241, T237};
  assign T237 = T239 ? T238 : 44'h0;
  assign T238 = ex_reg_pc;
  assign T239 = ex_reg_sel_alu1 == 2'h2;
  assign T240 = T5 ? io_ctrl_sel_alu1 : ex_reg_sel_alu1;
  assign T241 = T242 ? 20'hfffff : 20'h0;
  assign T242 = T237[6'h2b:6'h2b];
  assign T243 = ex_rs_0;
  assign T244 = ex_reg_sel_alu1 == 2'h1;
  assign T245 = ex_op2;
  assign ex_op2 = T316 ? T315 : T246;
  assign T246 = {T313, T247};
  assign T247 = T312 ? ex_imm : T248;
  assign T248 = {T252, T249};
  assign T249 = T250 ? 4'h4 : 4'h0;
  assign T250 = ex_reg_sel_alu2 == 3'h1;
  assign T251 = T5 ? io_ctrl_sel_alu2 : ex_reg_sel_alu2;
  assign T252 = T253 ? 28'hfffffff : 28'h0;
  assign T253 = T249[2'h3:2'h3];
  assign ex_imm = T254;
  assign T254 = {T298, T255};
  assign T255 = {T278, T256};
  assign T256 = {T267, T257};
  assign T257 = T266 ? T265 : T258;
  assign T258 = T264 ? T263 : T259;
  assign T259 = T261 ? T260 : 1'h0;
  assign T260 = ex_reg_inst[4'hf:4'hf];
  assign T261 = ex_reg_sel_imm == 3'h5;
  assign T262 = T5 ? io_ctrl_sel_imm : ex_reg_sel_imm;
  assign T263 = ex_reg_inst[5'h14:5'h14];
  assign T264 = ex_reg_sel_imm == 3'h4;
  assign T265 = ex_reg_inst[3'h7:3'h7];
  assign T266 = ex_reg_sel_imm == 3'h0;
  assign T267 = T277 ? 4'h0 : T268;
  assign T268 = T274 ? T273 : T269;
  assign T269 = T272 ? T271 : T270;
  assign T270 = ex_reg_inst[5'h18:5'h15];
  assign T271 = ex_reg_inst[5'h13:5'h10];
  assign T272 = ex_reg_sel_imm == 3'h5;
  assign T273 = ex_reg_inst[4'hb:4'h8];
  assign T274 = T276 | T275;
  assign T275 = ex_reg_sel_imm == 3'h1;
  assign T276 = ex_reg_sel_imm == 3'h0;
  assign T277 = ex_reg_sel_imm == 3'h2;
  assign T278 = {T284, T279};
  assign T279 = T281 ? 6'h0 : T280;
  assign T280 = ex_reg_inst[5'h1e:5'h19];
  assign T281 = T283 | T282;
  assign T282 = ex_reg_sel_imm == 3'h5;
  assign T283 = ex_reg_sel_imm == 3'h2;
  assign T284 = T295 ? 1'h0 : T285;
  assign T285 = T294 ? T292 : T286;
  assign T286 = T291 ? T289 : T287;
  assign T287 = T288;
  assign T288 = ex_reg_inst[5'h1f:5'h1f];
  assign T289 = T290;
  assign T290 = ex_reg_inst[3'h7:3'h7];
  assign T291 = ex_reg_sel_imm == 3'h1;
  assign T292 = T293;
  assign T293 = ex_reg_inst[5'h14:5'h14];
  assign T294 = ex_reg_sel_imm == 3'h3;
  assign T295 = T297 | T296;
  assign T296 = ex_reg_sel_imm == 3'h5;
  assign T297 = ex_reg_sel_imm == 3'h2;
  assign T298 = {T287, T299};
  assign T299 = {T307, T300};
  assign T300 = T304 ? T303 : T301;
  assign T301 = T302;
  assign T302 = ex_reg_inst[5'h13:4'hc];
  assign T303 = T287 ? 8'hff : 8'h0;
  assign T304 = T306 & T305;
  assign T305 = ex_reg_sel_imm != 3'h3;
  assign T306 = ex_reg_sel_imm != 3'h2;
  assign T307 = T311 ? T309 : T308;
  assign T308 = T287 ? 11'h7ff : 11'h0;
  assign T309 = T310;
  assign T310 = ex_reg_inst[5'h1e:5'h14];
  assign T311 = ex_reg_sel_imm == 3'h2;
  assign T312 = ex_reg_sel_alu2 == 3'h3;
  assign T313 = T314 ? 32'hffffffff : 32'h0;
  assign T314 = T247[5'h1f:5'h1f];
  assign T315 = ex_rs_1;
  assign T316 = ex_reg_sel_alu2 == 3'h2;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T135 = io_ctrl_mem_rocc_val ? mem_reg_rs2 : wb_reg_rs2;
  assign T136 = io_ctrl_ex_rs2_val ? ex_rs_1 : mem_reg_rs2;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_inst_opcode = T137;
  assign T137 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T138;
  assign T138 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T139;
  assign T139 = wb_reg_inst[4'hc:4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T140;
  assign T140 = wb_reg_inst[4'hd:4'hd];
  assign io_rocc_cmd_bits_inst_xd = T141;
  assign T141 = wb_reg_inst[4'he:4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T142;
  assign T142 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T143;
  assign T143 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T144;
  assign T144 = wb_reg_inst[5'h1f:5'h19];
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data;
  assign io_fpu_dmem_resp_tag = T211;
  assign T211 = dmem_resp_waddr[3'h4:1'h0];
  assign dmem_resp_waddr = T145 >> 1'h1;
  assign T145 = io_dmem_resp_bits_tag;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_val = T146;
  assign T146 = dmem_resp_valid & dmem_resp_fpu;
  assign dmem_resp_fpu = T147;
  assign T147 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign io_fpu_fcsr_rm = pcr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data;
  assign io_imem_btb_update_bits_returnAddr = T212;
  assign T212 = mem_int_wdata[6'h2a:1'h0];
  assign io_imem_btb_update_bits_target = T213;
  assign T213 = io_imem_req_bits_pc[6'h2a:1'h0];
  assign io_imem_btb_update_bits_pc = T214;
  assign T214 = mem_reg_pc[6'h2a:1'h0];
  assign io_imem_req_bits_pc = T215;
  assign T215 = T148[6'h2b:1'h0];
  assign T148 = T149;
  assign T149 = T167 ? mem_npc : T216;
  assign T216 = {1'h0, T150};
  assign T150 = T151 ? pcr_io_evec : wb_reg_pc;
  assign T151 = io_ctrl_sel_pc == 3'h3;
  assign mem_npc = io_ctrl_mem_jalr ? T217 : mem_br_target;
  assign T217 = {1'h0, T152};
  assign T152 = {T154, T153};
  assign T153 = mem_reg_wdata[6'h2a:1'h0];
  assign T154 = T164 ? T163 : T155;
  assign T155 = T159 ? T158 : T156;
  assign T156 = T157[1'h0:1'h0];
  assign T157 = mem_reg_wdata[6'h2b:6'h2a];
  assign T158 = T157 == 2'h3;
  assign T159 = T162 | T160;
  assign T160 = T161 == 22'h3ffffe;
  assign T161 = mem_reg_wdata >> 6'h2a;
  assign T162 = T161 == 22'h3fffff;
  assign T163 = T157 != 2'h0;
  assign T164 = T166 | T165;
  assign T165 = T161 == 22'h1;
  assign T166 = T161 == 22'h0;
  assign T167 = io_ctrl_sel_pc == 3'h1;
  assign io_ptw_status_s = pcr_io_status_s;
  assign io_ptw_status_ps = pcr_io_status_ps;
  assign io_ptw_status_ei = pcr_io_status_ei;
  assign io_ptw_status_pei = pcr_io_status_pei;
  assign io_ptw_status_ef = pcr_io_status_ef;
  assign io_ptw_status_u64 = pcr_io_status_u64;
  assign io_ptw_status_s64 = pcr_io_status_s64;
  assign io_ptw_status_vm = pcr_io_status_vm;
  assign io_ptw_status_er = pcr_io_status_er;
  assign io_ptw_status_zero = pcr_io_status_zero;
  assign io_ptw_status_im = pcr_io_status_im;
  assign io_ptw_status_ip = pcr_io_status_ip;
  assign io_ptw_sret = io_ctrl_sret;
  assign io_ptw_invalidate = pcr_io_fatc;
  assign io_ptw_ptbr = pcr_io_ptbr;
  assign io_dmem_req_bits_tag = T218;
  assign T218 = {2'h0, T168};
  assign T168 = {io_ctrl_ex_waddr, io_ctrl_ex_fp_val};
  assign io_dmem_req_bits_data = T169;
  assign T169 = io_ctrl_mem_fp_val ? io_fpu_store_data : mem_reg_rs2;
  assign io_dmem_req_bits_addr = T170;
  assign T170 = T171;
  assign T171 = {T173, T172};
  assign T172 = alu_io_adder_out[6'h2a:1'h0];
  assign T173 = T183 ? T182 : T174;
  assign T174 = T178 ? T177 : T175;
  assign T175 = T176[1'h0:1'h0];
  assign T176 = alu_io_adder_out[6'h2b:6'h2a];
  assign T177 = T176 == 2'h3;
  assign T178 = T181 | T179;
  assign T179 = T180 == 22'h3ffffe;
  assign T180 = ex_rs_0 >> 6'h2a;
  assign T181 = T180 == 22'h3fffff;
  assign T182 = T176 != 2'h0;
  assign T183 = T185 | T184;
  assign T184 = T180 == 22'h1;
  assign T185 = T180 == 22'h0;
  assign io_ctrl_csr_replay = pcr_io_replay;
  assign io_ctrl_fp_sboard_clra = T219;
  assign T219 = dmem_resp_waddr[3'h4:1'h0];
  assign io_ctrl_fp_sboard_clr = T186;
  assign T186 = dmem_resp_replay & dmem_resp_fpu;
  assign io_ctrl_status_s = pcr_io_status_s;
  assign io_ctrl_status_ps = pcr_io_status_ps;
  assign io_ctrl_status_ei = pcr_io_status_ei;
  assign io_ctrl_status_pei = pcr_io_status_pei;
  assign io_ctrl_status_ef = pcr_io_status_ef;
  assign io_ctrl_status_u64 = pcr_io_status_u64;
  assign io_ctrl_status_s64 = pcr_io_status_s64;
  assign io_ctrl_status_vm = pcr_io_status_vm;
  assign io_ctrl_status_er = pcr_io_status_er;
  assign io_ctrl_status_zero = pcr_io_status_zero;
  assign io_ctrl_status_im = pcr_io_status_im;
  assign io_ctrl_status_ip = pcr_io_status_ip;
  assign io_ctrl_wb_waddr = T187;
  assign T187 = wb_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_waddr = T188;
  assign T188 = mem_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_rs1_ra = T189;
  assign T189 = T190 == 5'h1;
  assign T190 = mem_reg_inst[5'h13:4'hf];
  assign io_ctrl_ex_waddr = T191;
  assign T191 = ex_reg_inst[4'hb:3'h7];
  assign io_ctrl_ll_waddr = T220;
  assign T220 = T192[3'h4:1'h0];
  assign T192 = T193 ? dmem_resp_waddr : T221;
  assign T221 = {2'h0, div_io_resp_bits_tag};
  assign io_ctrl_ll_wen = T194;
  assign T194 = T193 ? 1'h1 : T195;
  assign T195 = T232 & div_io_resp_valid;
  assign io_ctrl_div_mul_rdy = div_io_req_ready;
  assign io_ctrl_mem_misprediction = T196;
  assign T196 = T198 | T197;
  assign T197 = io_ctrl_ex_valid ^ 1'h1;
  assign T198 = mem_npc != T222;
  assign T222 = {1'h0, ex_reg_pc};
  assign io_ctrl_mem_br_taken = T199;
  assign T199 = mem_reg_wdata[1'h0:1'h0];
  assign io_ctrl_inst = io_imem_resp_bits_data;
  assign io_host_debug_stats_pcr = pcr_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = pcr_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = pcr_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = pcr_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = pcr_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = pcr_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = pcr_io_host_pcr_req_ready;
  ALU alu(
       .io_dw( ex_reg_ctrl_fn_dw ),
       .io_fn( ex_reg_ctrl_fn_alu ),
       .io_in2( T245 ),
       .io_in1( ex_op1 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( io_ctrl_div_mul_val ),
       .io_req_bits_fn( ex_reg_ctrl_fn_alu ),
       .io_req_bits_dw( ex_reg_ctrl_fn_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( io_ctrl_ex_waddr ),
       .io_kill( io_ctrl_div_mul_kill ),
       .io_resp_ready( T232 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );
  CSRFile pcr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( pcr_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( pcr_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( pcr_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( pcr_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( pcr_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( pcr_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( pcr_io_host_debug_stats_pcr ),
       .io_rw_addr( T231 ),
       .io_rw_cmd( T230 ),
       .io_rw_rdata( pcr_io_rw_rdata ),
       .io_rw_wdata( T223 ),
       .io_status_ip( pcr_io_status_ip ),
       .io_status_im( pcr_io_status_im ),
       .io_status_zero( pcr_io_status_zero ),
       .io_status_er( pcr_io_status_er ),
       .io_status_vm( pcr_io_status_vm ),
       .io_status_s64( pcr_io_status_s64 ),
       .io_status_u64( pcr_io_status_u64 ),
       .io_status_ef( pcr_io_status_ef ),
       .io_status_pei( pcr_io_status_pei ),
       .io_status_ei( pcr_io_status_ei ),
       .io_status_ps( pcr_io_status_ps ),
       .io_status_s( pcr_io_status_s ),
       .io_ptbr( pcr_io_ptbr ),
       .io_evec( pcr_io_evec ),
       .io_exception( io_ctrl_exception ),
       .io_retire( io_ctrl_retire ),
       .io_uarch_counters_15( 1'h0 ),
       .io_uarch_counters_14( 1'h0 ),
       .io_uarch_counters_13( 1'h0 ),
       .io_uarch_counters_12( 1'h0 ),
       .io_uarch_counters_11( 1'h0 ),
       .io_uarch_counters_10( 1'h0 ),
       .io_uarch_counters_9( 1'h0 ),
       .io_uarch_counters_8( 1'h0 ),
       .io_uarch_counters_7( 1'h0 ),
       .io_uarch_counters_6( 1'h0 ),
       .io_uarch_counters_5( 1'h0 ),
       .io_uarch_counters_4( 1'h0 ),
       .io_uarch_counters_3( 1'h0 ),
       .io_uarch_counters_2( 1'h0 ),
       .io_uarch_counters_1( 1'h0 ),
       .io_uarch_counters_0( 1'h0 ),
       .io_cause( io_ctrl_cause ),
       .io_badvaddr_wen( io_ctrl_badvaddr_wen ),
       .io_pc( wb_reg_pc ),
       .io_sret( io_ctrl_sret ),
       .io_fatc( pcr_io_fatc ),
       .io_replay( pcr_io_replay ),
       .io_time( pcr_io_time ),
       .io_fcsr_rm( pcr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );

  always @(posedge clk) begin
    if(T7) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T6) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data;
    end
    ex_reg_kill <= io_ctrl_killd;
    mem_reg_kill <= ex_reg_kill;
    R10 <= R11;
    if(ex_reg_rs_bypass_1) begin
      R11 <= T85;
    end else begin
      R11 <= T12;
    end
    if(T80) begin
      ex_reg_rs_lsb_1 <= io_ctrl_bypass_src_1;
    end else if(T79) begin
      ex_reg_rs_lsb_1 <= T15;
    end
    if (T20)
      T18[T25] <= wb_wdata;
    if(T7) begin
      wb_reg_wdata <= T32;
    end
    if(T6) begin
      mem_reg_wdata <= alu_io_out;
    end
    if(T6) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T83) begin
      ex_reg_rs_msb_1 <= T82;
    end
    if(T5) begin
      ex_reg_rs_bypass_1 <= io_ctrl_bypass_1;
    end
    R96 <= R97;
    if(ex_reg_rs_bypass_0) begin
      R97 <= T114;
    end else begin
      R97 <= T98;
    end
    if(T109) begin
      ex_reg_rs_lsb_0 <= io_ctrl_bypass_src_0;
    end else if(T108) begin
      ex_reg_rs_lsb_0 <= T101;
    end
    if(T112) begin
      ex_reg_rs_msb_0 <= T111;
    end
    if(T5) begin
      ex_reg_rs_bypass_0 <= io_ctrl_bypass_0;
    end
    if(T7) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if(T5) begin
      ex_reg_ctrl_fn_dw <= T234;
    end
    if(T5) begin
      ex_reg_ctrl_fn_alu <= io_ctrl_fn_alu;
    end
    if(T5) begin
      ex_reg_sel_alu1 <= io_ctrl_sel_alu1;
    end
    if(T5) begin
      ex_reg_sel_alu2 <= io_ctrl_sel_alu2;
    end
    if(T5) begin
      ex_reg_sel_imm <= io_ctrl_sel_imm;
    end
    if(io_ctrl_mem_rocc_val) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(io_ctrl_ex_rs2_val) begin
      mem_reg_rs2 <= ex_rs_1;
    end
`ifndef SYNTHESIS
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T133, T131, T130, T128, T126, T125, T124, T122, T95, T93, T9, T8, T1);
`endif
  end
endmodule

module Core(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    output io_imem_req_valid,
    output[43:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_index,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[2:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[3:0] io_imem_btb_update_bits_prediction_bits_bht_index,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_incorrectTarget,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    output[43:0] io_dmem_req_bits_addr,
    output[63:0] io_dmem_req_bits_data,
    output[7:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire[2:0] ctrl_io_dpath_sel_pc;
  wire ctrl_io_dpath_killd;
  wire ctrl_io_dpath_ren_1;
  wire ctrl_io_dpath_ren_0;
  wire[2:0] ctrl_io_dpath_sel_alu2;
  wire[1:0] ctrl_io_dpath_sel_alu1;
  wire[2:0] ctrl_io_dpath_sel_imm;
  wire ctrl_io_dpath_fn_dw;
  wire[3:0] ctrl_io_dpath_fn_alu;
  wire ctrl_io_dpath_div_mul_val;
  wire ctrl_io_dpath_div_mul_kill;
  wire[2:0] ctrl_io_dpath_csr;
  wire ctrl_io_dpath_sret;
  wire ctrl_io_dpath_mem_load;
  wire ctrl_io_dpath_wb_load;
  wire ctrl_io_dpath_ex_fp_val;
  wire ctrl_io_dpath_mem_fp_val;
  wire ctrl_io_dpath_ex_wen;
  wire ctrl_io_dpath_ex_valid;
  wire ctrl_io_dpath_mem_jalr;
  wire ctrl_io_dpath_mem_branch;
  wire ctrl_io_dpath_mem_wen;
  wire ctrl_io_dpath_wb_wen;
  wire[2:0] ctrl_io_dpath_ex_mem_type;
  wire ctrl_io_dpath_ex_rs2_val;
  wire ctrl_io_dpath_ex_rocc_val;
  wire ctrl_io_dpath_mem_rocc_val;
  wire ctrl_io_dpath_bypass_1;
  wire ctrl_io_dpath_bypass_0;
  wire[1:0] ctrl_io_dpath_bypass_src_1;
  wire[1:0] ctrl_io_dpath_bypass_src_0;
  wire ctrl_io_dpath_ll_ready;
  wire ctrl_io_dpath_retire;
  wire ctrl_io_dpath_exception;
  wire[63:0] ctrl_io_dpath_cause;
  wire ctrl_io_dpath_badvaddr_wen;
  wire ctrl_io_imem_req_valid;
  wire ctrl_io_imem_resp_ready;
  wire ctrl_io_imem_btb_update_valid;
  wire ctrl_io_imem_btb_update_bits_prediction_valid;
  wire ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  wire[42:0] ctrl_io_imem_btb_update_bits_prediction_bits_target;
  wire[2:0] ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  wire[3:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_index;
  wire[1:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire ctrl_io_imem_btb_update_bits_taken;
  wire ctrl_io_imem_btb_update_bits_isJump;
  wire ctrl_io_imem_btb_update_bits_isCall;
  wire ctrl_io_imem_btb_update_bits_isReturn;
  wire ctrl_io_imem_btb_update_bits_incorrectTarget;
  wire ctrl_io_imem_invalidate;
  wire ctrl_io_dmem_req_valid;
  wire ctrl_io_dmem_req_bits_kill;
  wire[2:0] ctrl_io_dmem_req_bits_typ;
  wire ctrl_io_dmem_req_bits_phys;
  wire[4:0] ctrl_io_dmem_req_bits_cmd;
  wire ctrl_io_rocc_cmd_valid;
  wire ctrl_io_rocc_s;
  wire ctrl_io_rocc_exception;
  wire dpath_io_host_pcr_req_ready;
  wire dpath_io_host_pcr_rep_valid;
  wire[63:0] dpath_io_host_pcr_rep_bits;
  wire dpath_io_host_ipi_req_valid;
  wire dpath_io_host_ipi_req_bits;
  wire dpath_io_host_ipi_rep_ready;
  wire dpath_io_host_debug_stats_pcr;
  wire[31:0] dpath_io_ctrl_inst;
  wire dpath_io_ctrl_mem_br_taken;
  wire dpath_io_ctrl_mem_misprediction;
  wire dpath_io_ctrl_div_mul_rdy;
  wire dpath_io_ctrl_ll_wen;
  wire[4:0] dpath_io_ctrl_ll_waddr;
  wire[4:0] dpath_io_ctrl_ex_waddr;
  wire dpath_io_ctrl_mem_rs1_ra;
  wire[4:0] dpath_io_ctrl_mem_waddr;
  wire[4:0] dpath_io_ctrl_wb_waddr;
  wire[7:0] dpath_io_ctrl_status_ip;
  wire[7:0] dpath_io_ctrl_status_im;
  wire[6:0] dpath_io_ctrl_status_zero;
  wire dpath_io_ctrl_status_er;
  wire dpath_io_ctrl_status_vm;
  wire dpath_io_ctrl_status_s64;
  wire dpath_io_ctrl_status_u64;
  wire dpath_io_ctrl_status_ef;
  wire dpath_io_ctrl_status_pei;
  wire dpath_io_ctrl_status_ei;
  wire dpath_io_ctrl_status_ps;
  wire dpath_io_ctrl_status_s;
  wire dpath_io_ctrl_fp_sboard_clr;
  wire[4:0] dpath_io_ctrl_fp_sboard_clra;
  wire dpath_io_ctrl_csr_replay;
  wire[43:0] dpath_io_dmem_req_bits_addr;
  wire[63:0] dpath_io_dmem_req_bits_data;
  wire[7:0] dpath_io_dmem_req_bits_tag;
  wire[31:0] dpath_io_ptw_ptbr;
  wire dpath_io_ptw_invalidate;
  wire dpath_io_ptw_sret;
  wire[7:0] dpath_io_ptw_status_ip;
  wire[7:0] dpath_io_ptw_status_im;
  wire[6:0] dpath_io_ptw_status_zero;
  wire dpath_io_ptw_status_er;
  wire dpath_io_ptw_status_vm;
  wire dpath_io_ptw_status_s64;
  wire dpath_io_ptw_status_u64;
  wire dpath_io_ptw_status_ef;
  wire dpath_io_ptw_status_pei;
  wire dpath_io_ptw_status_ei;
  wire dpath_io_ptw_status_ps;
  wire dpath_io_ptw_status_s;
  wire[43:0] dpath_io_imem_req_bits_pc;
  wire[42:0] dpath_io_imem_btb_update_bits_pc;
  wire[42:0] dpath_io_imem_btb_update_bits_target;
  wire[42:0] dpath_io_imem_btb_update_bits_returnAddr;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_funct;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs2;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs1;
  wire dpath_io_rocc_cmd_bits_inst_xd;
  wire dpath_io_rocc_cmd_bits_inst_xs1;
  wire dpath_io_rocc_cmd_bits_inst_xs2;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rd;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_opcode;
  wire[63:0] dpath_io_rocc_cmd_bits_rs1;
  wire[63:0] dpath_io_rocc_cmd_bits_rs2;


  assign io_rocc_exception = ctrl_io_rocc_exception;
  assign io_rocc_s = ctrl_io_rocc_s;
  assign io_rocc_cmd_bits_rs2 = dpath_io_rocc_cmd_bits_rs2;
  assign io_rocc_cmd_bits_rs1 = dpath_io_rocc_cmd_bits_rs1;
  assign io_rocc_cmd_bits_inst_opcode = dpath_io_rocc_cmd_bits_inst_opcode;
  assign io_rocc_cmd_bits_inst_rd = dpath_io_rocc_cmd_bits_inst_rd;
  assign io_rocc_cmd_bits_inst_xs2 = dpath_io_rocc_cmd_bits_inst_xs2;
  assign io_rocc_cmd_bits_inst_xs1 = dpath_io_rocc_cmd_bits_inst_xs1;
  assign io_rocc_cmd_bits_inst_xd = dpath_io_rocc_cmd_bits_inst_xd;
  assign io_rocc_cmd_bits_inst_rs1 = dpath_io_rocc_cmd_bits_inst_rs1;
  assign io_rocc_cmd_bits_inst_rs2 = dpath_io_rocc_cmd_bits_inst_rs2;
  assign io_rocc_cmd_bits_inst_funct = dpath_io_rocc_cmd_bits_inst_funct;
  assign io_rocc_cmd_valid = ctrl_io_rocc_cmd_valid;
  assign io_ptw_status_s = dpath_io_ptw_status_s;
  assign io_ptw_status_ps = dpath_io_ptw_status_ps;
  assign io_ptw_status_ei = dpath_io_ptw_status_ei;
  assign io_ptw_status_pei = dpath_io_ptw_status_pei;
  assign io_ptw_status_ef = dpath_io_ptw_status_ef;
  assign io_ptw_status_u64 = dpath_io_ptw_status_u64;
  assign io_ptw_status_s64 = dpath_io_ptw_status_s64;
  assign io_ptw_status_vm = dpath_io_ptw_status_vm;
  assign io_ptw_status_er = dpath_io_ptw_status_er;
  assign io_ptw_status_zero = dpath_io_ptw_status_zero;
  assign io_ptw_status_im = dpath_io_ptw_status_im;
  assign io_ptw_status_ip = dpath_io_ptw_status_ip;
  assign io_ptw_sret = dpath_io_ptw_sret;
  assign io_ptw_invalidate = dpath_io_ptw_invalidate;
  assign io_ptw_ptbr = dpath_io_ptw_ptbr;
  assign io_dmem_req_bits_cmd = ctrl_io_dmem_req_bits_cmd;
  assign io_dmem_req_bits_tag = dpath_io_dmem_req_bits_tag;
  assign io_dmem_req_bits_data = dpath_io_dmem_req_bits_data;
  assign io_dmem_req_bits_addr = dpath_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_phys = ctrl_io_dmem_req_bits_phys;
  assign io_dmem_req_bits_typ = ctrl_io_dmem_req_bits_typ;
  assign io_dmem_req_bits_kill = ctrl_io_dmem_req_bits_kill;
  assign io_dmem_req_valid = ctrl_io_dmem_req_valid;
  assign io_imem_invalidate = ctrl_io_imem_invalidate;
  assign io_imem_btb_update_bits_incorrectTarget = ctrl_io_imem_btb_update_bits_incorrectTarget;
  assign io_imem_btb_update_bits_isReturn = ctrl_io_imem_btb_update_bits_isReturn;
  assign io_imem_btb_update_bits_isCall = ctrl_io_imem_btb_update_bits_isCall;
  assign io_imem_btb_update_bits_isJump = ctrl_io_imem_btb_update_bits_isJump;
  assign io_imem_btb_update_bits_taken = ctrl_io_imem_btb_update_bits_taken;
  assign io_imem_btb_update_bits_returnAddr = dpath_io_imem_btb_update_bits_returnAddr;
  assign io_imem_btb_update_bits_target = dpath_io_imem_btb_update_bits_target;
  assign io_imem_btb_update_bits_pc = dpath_io_imem_btb_update_bits_pc;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_btb_update_bits_prediction_bits_bht_index = ctrl_io_imem_btb_update_bits_prediction_bits_bht_index;
  assign io_imem_btb_update_bits_prediction_bits_entry = ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = ctrl_io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_btb_update_bits_prediction_valid = ctrl_io_imem_btb_update_bits_prediction_valid;
  assign io_imem_btb_update_valid = ctrl_io_imem_btb_update_valid;
  assign io_imem_resp_ready = ctrl_io_imem_resp_ready;
  assign io_imem_req_bits_pc = dpath_io_imem_req_bits_pc;
  assign io_imem_req_valid = ctrl_io_imem_req_valid;
  assign io_host_debug_stats_pcr = dpath_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = dpath_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = dpath_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = dpath_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = dpath_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = dpath_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = dpath_io_host_pcr_req_ready;
  Control ctrl(.clk(clk), .reset(reset),
       .io_dpath_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_dpath_killd( ctrl_io_dpath_killd ),
       .io_dpath_ren_1( ctrl_io_dpath_ren_1 ),
       .io_dpath_ren_0( ctrl_io_dpath_ren_0 ),
       .io_dpath_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_dpath_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_dpath_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_dpath_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_dpath_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_dpath_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_dpath_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_dpath_div_val(  )
       //.io_dpath_div_kill(  )
       .io_dpath_csr( ctrl_io_dpath_csr ),
       .io_dpath_sret( ctrl_io_dpath_sret ),
       .io_dpath_mem_load( ctrl_io_dpath_mem_load ),
       .io_dpath_wb_load( ctrl_io_dpath_wb_load ),
       .io_dpath_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_dpath_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_dpath_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_dpath_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_dpath_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_dpath_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_dpath_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_dpath_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_dpath_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_dpath_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_dpath_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_dpath_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_dpath_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_dpath_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_dpath_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_dpath_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_dpath_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_dpath_retire( ctrl_io_dpath_retire ),
       .io_dpath_exception( ctrl_io_dpath_exception ),
       .io_dpath_cause( ctrl_io_dpath_cause ),
       .io_dpath_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_dpath_inst( dpath_io_ctrl_inst ),
       //.io_dpath_jalr_eq(  )
       .io_dpath_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_dpath_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_dpath_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_dpath_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_dpath_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_dpath_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_dpath_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_dpath_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_dpath_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_dpath_status_ip( dpath_io_ctrl_status_ip ),
       .io_dpath_status_im( dpath_io_ctrl_status_im ),
       .io_dpath_status_zero( dpath_io_ctrl_status_zero ),
       .io_dpath_status_er( dpath_io_ctrl_status_er ),
       .io_dpath_status_vm( dpath_io_ctrl_status_vm ),
       .io_dpath_status_s64( dpath_io_ctrl_status_s64 ),
       .io_dpath_status_u64( dpath_io_ctrl_status_u64 ),
       .io_dpath_status_ef( dpath_io_ctrl_status_ef ),
       .io_dpath_status_pei( dpath_io_ctrl_status_pei ),
       .io_dpath_status_ei( dpath_io_ctrl_status_ei ),
       .io_dpath_status_ps( dpath_io_ctrl_status_ps ),
       .io_dpath_status_s( dpath_io_ctrl_status_s ),
       .io_dpath_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_dpath_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_dpath_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_imem_req_valid( ctrl_io_imem_req_valid ),
       //.io_imem_req_bits_pc(  )
       .io_imem_resp_ready( ctrl_io_imem_resp_ready ),
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_index( io_imem_btb_resp_bits_bht_index ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( ctrl_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( ctrl_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( ctrl_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( ctrl_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( ctrl_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_index( ctrl_io_imem_btb_update_bits_prediction_bits_bht_index ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( ctrl_io_imem_btb_update_bits_prediction_bits_bht_value ),
       //.io_imem_btb_update_bits_pc(  )
       //.io_imem_btb_update_bits_target(  )
       //.io_imem_btb_update_bits_returnAddr(  )
       .io_imem_btb_update_bits_taken( ctrl_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( ctrl_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( ctrl_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( ctrl_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_incorrectTarget( ctrl_io_imem_btb_update_bits_incorrectTarget ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( ctrl_io_imem_invalidate ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       .io_dmem_req_valid( ctrl_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( ctrl_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( ctrl_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( ctrl_io_dmem_req_bits_phys ),
       //.io_dmem_req_bits_addr(  )
       //.io_dmem_req_bits_data(  )
       //.io_dmem_req_bits_tag(  )
       .io_dmem_req_bits_cmd( ctrl_io_dmem_req_bits_cmd ),
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       //.io_fpu_valid(  )
       //.io_fpu_fcsr_rdy(  )
       //.io_fpu_nack_mem(  )
       //.io_fpu_illegal_rm(  )
       //.io_fpu_killx(  )
       //.io_fpu_killm(  )
       //.io_fpu_dec_cmd(  )
       //.io_fpu_dec_ldst(  )
       //.io_fpu_dec_wen(  )
       //.io_fpu_dec_ren1(  )
       //.io_fpu_dec_ren2(  )
       //.io_fpu_dec_ren3(  )
       //.io_fpu_dec_swap23(  )
       //.io_fpu_dec_single(  )
       //.io_fpu_dec_fromint(  )
       //.io_fpu_dec_toint(  )
       //.io_fpu_dec_fastpipe(  )
       //.io_fpu_dec_fma(  )
       //.io_fpu_dec_round(  )
       //.io_fpu_sboard_set(  )
       //.io_fpu_sboard_clr(  )
       //.io_fpu_sboard_clra(  )
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( ctrl_io_rocc_cmd_valid ),
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       .io_rocc_s( ctrl_io_rocc_s ),
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       .io_rocc_exception( ctrl_io_rocc_exception )
  );
  `ifndef SYNTHESIS
    assign ctrl.io_fpu_nack_mem = {1{$random}};
    assign ctrl.io_fpu_illegal_rm = {1{$random}};
    assign ctrl.io_fpu_dec_wen = {1{$random}};
    assign ctrl.io_fpu_dec_ren1 = {1{$random}};
    assign ctrl.io_fpu_dec_ren2 = {1{$random}};
    assign ctrl.io_fpu_dec_ren3 = {1{$random}};
  `endif
  Datapath dpath(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( dpath_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( dpath_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( dpath_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( dpath_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( dpath_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( dpath_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( dpath_io_host_debug_stats_pcr ),
       .io_ctrl_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_ctrl_killd( ctrl_io_dpath_killd ),
       .io_ctrl_ren_1( ctrl_io_dpath_ren_1 ),
       .io_ctrl_ren_0( ctrl_io_dpath_ren_0 ),
       .io_ctrl_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_ctrl_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_ctrl_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_ctrl_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_ctrl_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_ctrl_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_ctrl_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_ctrl_div_val(  )
       //.io_ctrl_div_kill(  )
       .io_ctrl_csr( ctrl_io_dpath_csr ),
       .io_ctrl_sret( ctrl_io_dpath_sret ),
       .io_ctrl_mem_load( ctrl_io_dpath_mem_load ),
       .io_ctrl_wb_load( ctrl_io_dpath_wb_load ),
       .io_ctrl_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_ctrl_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_ctrl_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_ctrl_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_ctrl_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_ctrl_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_ctrl_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_ctrl_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_ctrl_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_ctrl_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_ctrl_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_ctrl_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_ctrl_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_ctrl_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_ctrl_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_ctrl_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_ctrl_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_ctrl_retire( ctrl_io_dpath_retire ),
       .io_ctrl_exception( ctrl_io_dpath_exception ),
       .io_ctrl_cause( ctrl_io_dpath_cause ),
       .io_ctrl_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_ctrl_inst( dpath_io_ctrl_inst ),
       //.io_ctrl_jalr_eq(  )
       .io_ctrl_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_ctrl_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_ctrl_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_ctrl_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_ctrl_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_ctrl_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_ctrl_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_ctrl_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_ctrl_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_ctrl_status_ip( dpath_io_ctrl_status_ip ),
       .io_ctrl_status_im( dpath_io_ctrl_status_im ),
       .io_ctrl_status_zero( dpath_io_ctrl_status_zero ),
       .io_ctrl_status_er( dpath_io_ctrl_status_er ),
       .io_ctrl_status_vm( dpath_io_ctrl_status_vm ),
       .io_ctrl_status_s64( dpath_io_ctrl_status_s64 ),
       .io_ctrl_status_u64( dpath_io_ctrl_status_u64 ),
       .io_ctrl_status_ef( dpath_io_ctrl_status_ef ),
       .io_ctrl_status_pei( dpath_io_ctrl_status_pei ),
       .io_ctrl_status_ei( dpath_io_ctrl_status_ei ),
       .io_ctrl_status_ps( dpath_io_ctrl_status_ps ),
       .io_ctrl_status_s( dpath_io_ctrl_status_s ),
       .io_ctrl_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_ctrl_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_ctrl_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       //.io_dmem_req_valid(  )
       //.io_dmem_req_bits_kill(  )
       //.io_dmem_req_bits_typ(  )
       //.io_dmem_req_bits_phys(  )
       .io_dmem_req_bits_addr( dpath_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_data( dpath_io_dmem_req_bits_data ),
       .io_dmem_req_bits_tag( dpath_io_dmem_req_bits_tag ),
       //.io_dmem_req_bits_cmd(  )
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_ptw_ptbr( dpath_io_ptw_ptbr ),
       .io_ptw_invalidate( dpath_io_ptw_invalidate ),
       .io_ptw_sret( dpath_io_ptw_sret ),
       .io_ptw_status_ip( dpath_io_ptw_status_ip ),
       .io_ptw_status_im( dpath_io_ptw_status_im ),
       .io_ptw_status_zero( dpath_io_ptw_status_zero ),
       .io_ptw_status_er( dpath_io_ptw_status_er ),
       .io_ptw_status_vm( dpath_io_ptw_status_vm ),
       .io_ptw_status_s64( dpath_io_ptw_status_s64 ),
       .io_ptw_status_u64( dpath_io_ptw_status_u64 ),
       .io_ptw_status_ef( dpath_io_ptw_status_ef ),
       .io_ptw_status_pei( dpath_io_ptw_status_pei ),
       .io_ptw_status_ei( dpath_io_ptw_status_ei ),
       .io_ptw_status_ps( dpath_io_ptw_status_ps ),
       .io_ptw_status_s( dpath_io_ptw_status_s ),
       //.io_imem_req_valid(  )
       .io_imem_req_bits_pc( dpath_io_imem_req_bits_pc ),
       //.io_imem_resp_ready(  )
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_index( io_imem_btb_resp_bits_bht_index ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       //.io_imem_btb_update_valid(  )
       //.io_imem_btb_update_bits_prediction_valid(  )
       //.io_imem_btb_update_bits_prediction_bits_taken(  )
       //.io_imem_btb_update_bits_prediction_bits_target(  )
       //.io_imem_btb_update_bits_prediction_bits_entry(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_index(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_value(  )
       .io_imem_btb_update_bits_pc( dpath_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( dpath_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( dpath_io_imem_btb_update_bits_returnAddr ),
       //.io_imem_btb_update_bits_taken(  )
       //.io_imem_btb_update_bits_isJump(  )
       //.io_imem_btb_update_bits_isCall(  )
       //.io_imem_btb_update_bits_isReturn(  )
       //.io_imem_btb_update_bits_incorrectTarget(  )
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       //.io_imem_invalidate(  )
       //.io_fpu_inst(  )
       //.io_fpu_fromint_data(  )
       //.io_fpu_fcsr_rm(  )
       //.io_fpu_fcsr_flags_valid(  )
       //.io_fpu_fcsr_flags_bits(  )
       //.io_fpu_store_data(  )
       //.io_fpu_toint_data(  )
       //.io_fpu_dmem_resp_val(  )
       //.io_fpu_dmem_resp_type(  )
       //.io_fpu_dmem_resp_tag(  )
       //.io_fpu_dmem_resp_data(  )
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       .io_rocc_cmd_bits_inst_funct( dpath_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( dpath_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( dpath_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( dpath_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( dpath_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( dpath_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( dpath_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( dpath_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( dpath_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( dpath_io_rocc_cmd_bits_rs2 ),
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );
  `ifndef SYNTHESIS
    assign dpath.io_fpu_fcsr_flags_valid = {1{$random}};
    assign dpath.io_fpu_fcsr_flags_bits = {1{$random}};
    assign dpath.io_fpu_store_data = {2{$random}};
    assign dpath.io_fpu_toint_data = {2{$random}};
  `endif
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input  io_requestor_1_req_bits_kill,
    input [2:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_phys,
    input [43:0] io_requestor_1_req_bits_addr,
    input [63:0] io_requestor_1_req_bits_data,
    input [7:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output[2:0] io_requestor_1_resp_bits_typ,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data,
    output[63:0] io_requestor_1_resp_bits_data_subword,
    output[7:0] io_requestor_1_resp_bits_tag,
    output[3:0] io_requestor_1_resp_bits_cmd,
    output[43:0] io_requestor_1_resp_bits_addr,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[7:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    //input  io_requestor_1_ptw_req_ready
    //output io_requestor_1_ptw_req_valid
    //output[29:0] io_requestor_1_ptw_req_bits
    //input  io_requestor_1_ptw_resp_valid
    //input  io_requestor_1_ptw_resp_bits_error
    //input [18:0] io_requestor_1_ptw_resp_bits_ppn
    //input [5:0] io_requestor_1_ptw_resp_bits_perm
    //input [7:0] io_requestor_1_ptw_status_ip
    //input [7:0] io_requestor_1_ptw_status_im
    //input [6:0] io_requestor_1_ptw_status_zero
    //input  io_requestor_1_ptw_status_er
    //input  io_requestor_1_ptw_status_vm
    //input  io_requestor_1_ptw_status_s64
    //input  io_requestor_1_ptw_status_u64
    //input  io_requestor_1_ptw_status_ef
    //input  io_requestor_1_ptw_status_pei
    //input  io_requestor_1_ptw_status_ei
    //input  io_requestor_1_ptw_status_ps
    //input  io_requestor_1_ptw_status_s
    //input  io_requestor_1_ptw_invalidate
    //input  io_requestor_1_ptw_sret
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input  io_requestor_0_req_bits_kill,
    input [2:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_phys,
    input [43:0] io_requestor_0_req_bits_addr,
    input [63:0] io_requestor_0_req_bits_data,
    input [7:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output[2:0] io_requestor_0_resp_bits_typ,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data,
    output[63:0] io_requestor_0_resp_bits_data_subword,
    output[7:0] io_requestor_0_resp_bits_tag,
    output[3:0] io_requestor_0_resp_bits_cmd,
    output[43:0] io_requestor_0_resp_bits_addr,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[7:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_ptw_req_ready
    //output io_requestor_0_ptw_req_valid
    //output[29:0] io_requestor_0_ptw_req_bits
    //input  io_requestor_0_ptw_resp_valid
    //input  io_requestor_0_ptw_resp_bits_error
    //input [18:0] io_requestor_0_ptw_resp_bits_ppn
    //input [5:0] io_requestor_0_ptw_resp_bits_perm
    //input [7:0] io_requestor_0_ptw_status_ip
    //input [7:0] io_requestor_0_ptw_status_im
    //input [6:0] io_requestor_0_ptw_status_zero
    //input  io_requestor_0_ptw_status_er
    //input  io_requestor_0_ptw_status_vm
    //input  io_requestor_0_ptw_status_s64
    //input  io_requestor_0_ptw_status_u64
    //input  io_requestor_0_ptw_status_ef
    //input  io_requestor_0_ptw_status_pei
    //input  io_requestor_0_ptw_status_ei
    //input  io_requestor_0_ptw_status_ps
    //input  io_requestor_0_ptw_status_s
    //input  io_requestor_0_ptw_invalidate
    //input  io_requestor_0_ptw_sret
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    output[63:0] io_mem_req_bits_data,
    output[7:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    input  io_mem_resp_valid,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    input  io_mem_ptw_req_valid,
    input [29:0] io_mem_ptw_req_bits,
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered
);

  wire[4:0] T0;
  wire[7:0] T32;
  wire[8:0] T1;
  wire[8:0] T2;
  wire[8:0] T3;
  wire[63:0] T4;
  reg  r_valid_0;
  wire[43:0] T5;
  wire T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  wire[7:0] T33;
  wire[6:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire[7:0] T34;
  wire[6:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[7:0] T35;
  wire[6:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[7:0] T36;
  wire[6:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_valid_0 = {1{$random}};
  end
`endif

  assign io_mem_req_bits_cmd = T0;
  assign T0 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign io_mem_req_bits_tag = T32;
  assign T32 = T1[3'h7:1'h0];
  assign T1 = io_requestor_0_req_valid ? T3 : T2;
  assign T2 = {io_requestor_1_req_bits_tag, 1'h1};
  assign T3 = {io_requestor_0_req_bits_tag, 1'h0};
  assign io_mem_req_bits_data = T4;
  assign T4 = r_valid_0 ? io_requestor_0_req_bits_data : io_requestor_1_req_bits_data;
  assign io_mem_req_bits_addr = T5;
  assign T5 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign io_mem_req_bits_phys = T6;
  assign T6 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign io_mem_req_bits_typ = T7;
  assign T7 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign io_mem_req_bits_kill = T8;
  assign T8 = r_valid_0 ? io_requestor_0_req_bits_kill : io_requestor_1_req_bits_kill;
  assign io_mem_req_valid = T9;
  assign T9 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T33;
  assign T33 = {1'h0, T10};
  assign T10 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_0_replay_next_valid = T11;
  assign T11 = io_mem_replay_next_valid & T12;
  assign T12 = T13 == 1'h0;
  assign T13 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T34;
  assign T34 = {1'h0, T14};
  assign T14 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_0_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_replay = T15;
  assign T15 = io_mem_resp_bits_replay & T16;
  assign T16 = T17 == 1'h0;
  assign T17 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_0_resp_bits_nack = T18;
  assign T18 = io_mem_resp_bits_nack & T16;
  assign io_requestor_0_resp_valid = T19;
  assign T19 = io_mem_resp_valid & T16;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T35;
  assign T35 = {1'h0, T20};
  assign T20 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_1_replay_next_valid = T21;
  assign T21 = io_mem_replay_next_valid & T22;
  assign T22 = T23 == 1'h1;
  assign T23 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T36;
  assign T36 = {1'h0, T24};
  assign T24 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_1_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_replay = T25;
  assign T25 = io_mem_resp_bits_replay & T26;
  assign T26 = T27 == 1'h1;
  assign T27 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_1_resp_bits_nack = T28;
  assign T28 = io_mem_resp_bits_nack & T26;
  assign io_requestor_1_resp_valid = T29;
  assign T29 = io_mem_resp_valid & T26;
  assign io_requestor_1_req_ready = T30;
  assign T30 = io_requestor_0_req_ready & T31;
  assign T31 = io_requestor_0_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T36;
  wire T6;
  wire T7;
  wire[3:0] T8;
  wire T9;
  wire[2:0] T10;
  wire[5:0] T11;
  wire[2:0] T12;
  wire[511:0] T13;
  wire[1:0] T14;
  wire[25:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T36 = reset ? 1'h0 : T6;
  assign T6 = T7 ? T0 : R5;
  assign T7 = io_out_ready & io_out_valid;
  assign io_out_bits_payload_atomic_opcode = T8;
  assign T8 = T9 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T9 = T0;
  assign io_out_bits_payload_subword_addr = T10;
  assign T10 = T9 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign io_out_bits_payload_write_mask = T11;
  assign T11 = T9 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign io_out_bits_payload_a_type = T12;
  assign T12 = T9 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign io_out_bits_payload_data = T13;
  assign T13 = T9 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign io_out_bits_payload_client_xact_id = T14;
  assign T14 = T9 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign io_out_bits_payload_addr = T15;
  assign T15 = T9 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign io_out_bits_header_dst = T16;
  assign T16 = T9 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T17;
  assign T17 = T9 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T18;
  assign T18 = T9 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T19;
  assign T19 = T20 & io_out_ready;
  assign T20 = T27 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = T25 | T23;
  assign T23 = io_in_1_valid & T24;
  assign T24 = R5 < 1'h1;
  assign T25 = io_in_0_valid & T26;
  assign T26 = R5 < 1'h0;
  assign T27 = R5 < 1'h0;
  assign io_in_1_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = T33 | T30;
  assign T30 = T31 ^ 1'h1;
  assign T31 = T32 | io_in_0_valid;
  assign T32 = T25 | T23;
  assign T33 = T35 & T34;
  assign T34 = R5 < 1'h1;
  assign T35 = T25 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T7) begin
      R5 <= T0;
    end
  end
endmodule

module RRArbiter_2(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T30;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T30 = reset ? 1'h0 : T6;
  assign T6 = T7 ? T0 : R5;
  assign T7 = io_out_ready & io_out_valid;
  assign io_out_bits_payload_master_xact_id = T8;
  assign T8 = T9 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T9 = T0;
  assign io_out_bits_header_dst = T10;
  assign T10 = T9 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T11;
  assign T11 = T9 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T12;
  assign T12 = T9 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T13;
  assign T13 = T14 & io_out_ready;
  assign T14 = T21 | T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = T19 | T17;
  assign T17 = io_in_1_valid & T18;
  assign T18 = R5 < 1'h1;
  assign T19 = io_in_0_valid & T20;
  assign T20 = R5 < 1'h0;
  assign T21 = R5 < 1'h0;
  assign io_in_1_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = T27 | T24;
  assign T24 = T25 ^ 1'h1;
  assign T25 = T26 | io_in_0_valid;
  assign T26 = T19 | T17;
  assign T27 = T29 & T28;
  assign T28 = R5 < 1'h1;
  assign T29 = T19 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T7) begin
      R5 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatAppendsArbiterId(input clk, input reset,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [1:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_1_acquire_bits_payload_data,
    input [2:0] io_in_1_acquire_bits_payload_a_type,
    input [5:0] io_in_1_acquire_bits_payload_write_mask,
    input [2:0] io_in_1_acquire_bits_payload_subword_addr,
    input [3:0] io_in_1_acquire_bits_payload_atomic_opcode,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[511:0] io_in_1_grant_bits_payload_data,
    output[1:0] io_in_1_grant_bits_payload_client_xact_id,
    output[2:0] io_in_1_grant_bits_payload_master_xact_id,
    output[3:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input [2:0] io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [1:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_0_acquire_bits_payload_data,
    input [2:0] io_in_0_acquire_bits_payload_a_type,
    input [5:0] io_in_0_acquire_bits_payload_write_mask,
    input [2:0] io_in_0_acquire_bits_payload_subword_addr,
    input [3:0] io_in_0_acquire_bits_payload_atomic_opcode,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[511:0] io_in_0_grant_bits_payload_data,
    output[1:0] io_in_0_grant_bits_payload_client_xact_id,
    output[2:0] io_in_0_grant_bits_payload_master_xact_id,
    output[3:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input [2:0] io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[1:0] io_out_acquire_bits_payload_client_xact_id,
    output[511:0] io_out_acquire_bits_payload_data,
    output[2:0] io_out_acquire_bits_payload_a_type,
    output[5:0] io_out_acquire_bits_payload_write_mask,
    output[2:0] io_out_acquire_bits_payload_subword_addr,
    output[3:0] io_out_acquire_bits_payload_atomic_opcode,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [511:0] io_out_grant_bits_payload_data,
    input [1:0] io_out_grant_bits_payload_client_xact_id,
    input [2:0] io_out_grant_bits_payload_master_xact_id,
    input [3:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[2:0] io_out_finish_bits_payload_master_xact_id
);

  wire[1:0] T14;
  wire[2:0] T15;
  wire[1:0] T16;
  wire[2:0] T17;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[1:0] T12;
  wire T8;
  wire T9;
  wire[1:0] T13;
  wire T10;
  wire T11;
  wire RRArbiter_0_io_in_1_ready;
  wire RRArbiter_0_io_in_0_ready;
  wire RRArbiter_0_io_out_valid;
  wire[1:0] RRArbiter_0_io_out_bits_header_src;
  wire[1:0] RRArbiter_0_io_out_bits_header_dst;
  wire[25:0] RRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] RRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[511:0] RRArbiter_0_io_out_bits_payload_data;
  wire[2:0] RRArbiter_0_io_out_bits_payload_a_type;
  wire[5:0] RRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] RRArbiter_0_io_out_bits_payload_subword_addr;
  wire[3:0] RRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire RRArbiter_1_io_in_1_ready;
  wire RRArbiter_1_io_in_0_ready;
  wire RRArbiter_1_io_out_valid;
  wire[1:0] RRArbiter_1_io_out_bits_header_src;
  wire[1:0] RRArbiter_1_io_out_bits_header_dst;
  wire[2:0] RRArbiter_1_io_out_bits_payload_master_xact_id;


  assign T14 = T15[1'h1:1'h0];
  assign T15 = {io_in_0_acquire_bits_payload_client_xact_id, 1'h0};
  assign T16 = T17[1'h1:1'h0];
  assign T17 = {io_in_1_acquire_bits_payload_client_xact_id, 1'h1};
  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_1_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_1_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_1_io_out_valid;
  assign io_out_grant_ready = T0;
  assign T0 = T5 ? io_in_1_grant_ready : T1;
  assign T1 = T2 ? io_in_0_grant_ready : 1'h0;
  assign T2 = T3 == 1'h0;
  assign T3 = T4;
  assign T4 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign T5 = T6 == 1'h1;
  assign T6 = T7;
  assign T7 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_out_acquire_bits_payload_atomic_opcode = RRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_acquire_bits_payload_subword_addr = RRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_acquire_bits_payload_write_mask = RRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_data = RRArbiter_0_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_0_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_0_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_0_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_0_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_1_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = T12;
  assign T12 = {1'h0, T8};
  assign T8 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T9;
  assign T9 = T2 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_0_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_1_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = T13;
  assign T13 = {1'h0, T10};
  assign T10 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T11;
  assign T11 = T5 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_0_io_in_1_ready;
  RRArbiter_1 RRArbiter_0(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( T16 ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_acquire_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_acquire_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_acquire_bits_payload_atomic_opcode ),
       .io_in_0_ready( RRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( T14 ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_acquire_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_acquire_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_acquire_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( RRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( RRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( RRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( RRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  RRArbiter_2 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_1_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module Tile(input clk, input reset,
    input  io_tilelink_acquire_ready,
    output io_tilelink_acquire_valid,
    output[1:0] io_tilelink_acquire_bits_header_src,
    output[1:0] io_tilelink_acquire_bits_header_dst,
    output[25:0] io_tilelink_acquire_bits_payload_addr,
    output[1:0] io_tilelink_acquire_bits_payload_client_xact_id,
    output[511:0] io_tilelink_acquire_bits_payload_data,
    output[2:0] io_tilelink_acquire_bits_payload_a_type,
    output[5:0] io_tilelink_acquire_bits_payload_write_mask,
    output[2:0] io_tilelink_acquire_bits_payload_subword_addr,
    output[3:0] io_tilelink_acquire_bits_payload_atomic_opcode,
    output io_tilelink_grant_ready,
    input  io_tilelink_grant_valid,
    input [1:0] io_tilelink_grant_bits_header_src,
    input [1:0] io_tilelink_grant_bits_header_dst,
    input [511:0] io_tilelink_grant_bits_payload_data,
    input [1:0] io_tilelink_grant_bits_payload_client_xact_id,
    input [2:0] io_tilelink_grant_bits_payload_master_xact_id,
    input [3:0] io_tilelink_grant_bits_payload_g_type,
    input  io_tilelink_finish_ready,
    output io_tilelink_finish_valid,
    output[1:0] io_tilelink_finish_bits_header_src,
    output[1:0] io_tilelink_finish_bits_header_dst,
    output[2:0] io_tilelink_finish_bits_payload_master_xact_id,
    output io_tilelink_probe_ready,
    input  io_tilelink_probe_valid,
    input [1:0] io_tilelink_probe_bits_header_src,
    input [1:0] io_tilelink_probe_bits_header_dst,
    input [25:0] io_tilelink_probe_bits_payload_addr,
    input [2:0] io_tilelink_probe_bits_payload_master_xact_id,
    input [1:0] io_tilelink_probe_bits_payload_p_type,
    input  io_tilelink_release_ready,
    output io_tilelink_release_valid,
    output[1:0] io_tilelink_release_bits_header_src,
    output[1:0] io_tilelink_release_bits_header_dst,
    output[25:0] io_tilelink_release_bits_payload_addr,
    output[1:0] io_tilelink_release_bits_payload_client_xact_id,
    output[2:0] io_tilelink_release_bits_payload_master_xact_id,
    output[511:0] io_tilelink_release_bits_payload_data,
    output[2:0] io_tilelink_release_bits_payload_r_type,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr
);

  wire[1:0] T1;
  wire[2:0] T0;
  wire dcArb_io_requestor_1_req_ready;
  wire dcArb_io_requestor_1_resp_valid;
  wire dcArb_io_requestor_1_resp_bits_nack;
  wire dcArb_io_requestor_1_resp_bits_replay;
  wire[2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire dcArb_io_requestor_1_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data_subword;
  wire[7:0] dcArb_io_requestor_1_resp_bits_tag;
  wire[3:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire[43:0] dcArb_io_requestor_1_resp_bits_addr;
  wire[63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire dcArb_io_requestor_1_replay_next_valid;
  wire[7:0] dcArb_io_requestor_1_replay_next_bits;
  wire dcArb_io_requestor_1_xcpt_ma_ld;
  wire dcArb_io_requestor_1_xcpt_ma_st;
  wire dcArb_io_requestor_1_xcpt_pf_ld;
  wire dcArb_io_requestor_1_xcpt_pf_st;
  wire dcArb_io_requestor_1_ordered;
  wire dcArb_io_requestor_0_req_ready;
  wire dcArb_io_requestor_0_resp_valid;
  wire dcArb_io_requestor_0_resp_bits_nack;
  wire dcArb_io_requestor_0_resp_bits_replay;
  wire[2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire dcArb_io_requestor_0_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data_subword;
  wire[7:0] dcArb_io_requestor_0_resp_bits_tag;
  wire[3:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire[43:0] dcArb_io_requestor_0_resp_bits_addr;
  wire[63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire dcArb_io_requestor_0_replay_next_valid;
  wire[7:0] dcArb_io_requestor_0_replay_next_bits;
  wire dcArb_io_requestor_0_xcpt_ma_ld;
  wire dcArb_io_requestor_0_xcpt_ma_st;
  wire dcArb_io_requestor_0_xcpt_pf_ld;
  wire dcArb_io_requestor_0_xcpt_pf_st;
  wire dcArb_io_requestor_0_ordered;
  wire dcArb_io_mem_req_valid;
  wire dcArb_io_mem_req_bits_kill;
  wire[2:0] dcArb_io_mem_req_bits_typ;
  wire dcArb_io_mem_req_bits_phys;
  wire[43:0] dcArb_io_mem_req_bits_addr;
  wire[63:0] dcArb_io_mem_req_bits_data;
  wire[7:0] dcArb_io_mem_req_bits_tag;
  wire[4:0] dcArb_io_mem_req_bits_cmd;
  wire ptw_io_requestor_1_req_ready;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_resp_bits_error;
  wire[18:0] ptw_io_requestor_1_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_1_resp_bits_perm;
  wire[7:0] ptw_io_requestor_1_status_ip;
  wire[7:0] ptw_io_requestor_1_status_im;
  wire[6:0] ptw_io_requestor_1_status_zero;
  wire ptw_io_requestor_1_status_er;
  wire ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_s64;
  wire ptw_io_requestor_1_status_u64;
  wire ptw_io_requestor_1_status_ef;
  wire ptw_io_requestor_1_status_pei;
  wire ptw_io_requestor_1_status_ei;
  wire ptw_io_requestor_1_status_ps;
  wire ptw_io_requestor_1_status_s;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_1_sret;
  wire ptw_io_requestor_0_req_ready;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_resp_bits_error;
  wire[18:0] ptw_io_requestor_0_resp_bits_ppn;
  wire[5:0] ptw_io_requestor_0_resp_bits_perm;
  wire[7:0] ptw_io_requestor_0_status_ip;
  wire[7:0] ptw_io_requestor_0_status_im;
  wire[6:0] ptw_io_requestor_0_status_zero;
  wire ptw_io_requestor_0_status_er;
  wire ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_s64;
  wire ptw_io_requestor_0_status_u64;
  wire ptw_io_requestor_0_status_ef;
  wire ptw_io_requestor_0_status_pei;
  wire ptw_io_requestor_0_status_ei;
  wire ptw_io_requestor_0_status_ps;
  wire ptw_io_requestor_0_status_s;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_requestor_0_sret;
  wire ptw_io_mem_req_valid;
  wire ptw_io_mem_req_bits_kill;
  wire[2:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_phys;
  wire[43:0] ptw_io_mem_req_bits_addr;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire memArb_io_in_1_acquire_ready;
  wire memArb_io_in_1_grant_valid;
  wire[1:0] memArb_io_in_1_grant_bits_header_src;
  wire[1:0] memArb_io_in_1_grant_bits_header_dst;
  wire[511:0] memArb_io_in_1_grant_bits_payload_data;
  wire[1:0] memArb_io_in_1_grant_bits_payload_client_xact_id;
  wire[2:0] memArb_io_in_1_grant_bits_payload_master_xact_id;
  wire[3:0] memArb_io_in_1_grant_bits_payload_g_type;
  wire memArb_io_in_1_finish_ready;
  wire memArb_io_in_0_acquire_ready;
  wire memArb_io_in_0_grant_valid;
  wire[1:0] memArb_io_in_0_grant_bits_header_src;
  wire[1:0] memArb_io_in_0_grant_bits_header_dst;
  wire[511:0] memArb_io_in_0_grant_bits_payload_data;
  wire[1:0] memArb_io_in_0_grant_bits_payload_client_xact_id;
  wire[2:0] memArb_io_in_0_grant_bits_payload_master_xact_id;
  wire[3:0] memArb_io_in_0_grant_bits_payload_g_type;
  wire memArb_io_in_0_finish_ready;
  wire memArb_io_out_acquire_valid;
  wire[1:0] memArb_io_out_acquire_bits_header_src;
  wire[1:0] memArb_io_out_acquire_bits_header_dst;
  wire[25:0] memArb_io_out_acquire_bits_payload_addr;
  wire[1:0] memArb_io_out_acquire_bits_payload_client_xact_id;
  wire[511:0] memArb_io_out_acquire_bits_payload_data;
  wire[2:0] memArb_io_out_acquire_bits_payload_a_type;
  wire[5:0] memArb_io_out_acquire_bits_payload_write_mask;
  wire[2:0] memArb_io_out_acquire_bits_payload_subword_addr;
  wire[3:0] memArb_io_out_acquire_bits_payload_atomic_opcode;
  wire memArb_io_out_grant_ready;
  wire memArb_io_out_finish_valid;
  wire[1:0] memArb_io_out_finish_bits_header_src;
  wire[1:0] memArb_io_out_finish_bits_header_dst;
  wire[2:0] memArb_io_out_finish_bits_payload_master_xact_id;
  wire icache_io_cpu_resp_valid;
  wire[43:0] icache_io_cpu_resp_bits_pc;
  wire[31:0] icache_io_cpu_resp_bits_data;
  wire icache_io_cpu_resp_bits_xcpt_ma;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire[42:0] icache_io_cpu_btb_resp_bits_target;
  wire[2:0] icache_io_cpu_btb_resp_bits_entry;
  wire[3:0] icache_io_cpu_btb_resp_bits_bht_index;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire icache_io_cpu_ptw_req_valid;
  wire[29:0] icache_io_cpu_ptw_req_bits;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire[1:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire[2:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[5:0] icache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] icache_io_mem_acquire_bits_payload_subword_addr;
  wire[3:0] icache_io_mem_acquire_bits_payload_atomic_opcode;
  wire icache_io_mem_grant_ready;
  wire icache_io_mem_finish_valid;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[2:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire core_io_host_pcr_req_ready;
  wire core_io_host_pcr_rep_valid;
  wire[63:0] core_io_host_pcr_rep_bits;
  wire core_io_host_ipi_req_valid;
  wire core_io_host_ipi_req_bits;
  wire core_io_host_ipi_rep_ready;
  wire core_io_host_debug_stats_pcr;
  wire core_io_imem_req_valid;
  wire[43:0] core_io_imem_req_bits_pc;
  wire core_io_imem_resp_ready;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire[42:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire[2:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[3:0] core_io_imem_btb_update_bits_prediction_bits_bht_index;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[42:0] core_io_imem_btb_update_bits_pc;
  wire[42:0] core_io_imem_btb_update_bits_target;
  wire[42:0] core_io_imem_btb_update_bits_returnAddr;
  wire core_io_imem_btb_update_bits_taken;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_isCall;
  wire core_io_imem_btb_update_bits_isReturn;
  wire core_io_imem_btb_update_bits_incorrectTarget;
  wire core_io_imem_invalidate;
  wire core_io_dmem_req_valid;
  wire core_io_dmem_req_bits_kill;
  wire[2:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_phys;
  wire[43:0] core_io_dmem_req_bits_addr;
  wire[63:0] core_io_dmem_req_bits_data;
  wire[7:0] core_io_dmem_req_bits_tag;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[31:0] core_io_ptw_ptbr;
  wire core_io_ptw_invalidate;
  wire core_io_ptw_sret;
  wire[7:0] core_io_ptw_status_ip;
  wire[7:0] core_io_ptw_status_im;
  wire[6:0] core_io_ptw_status_zero;
  wire core_io_ptw_status_er;
  wire core_io_ptw_status_vm;
  wire core_io_ptw_status_s64;
  wire core_io_ptw_status_u64;
  wire core_io_ptw_status_ef;
  wire core_io_ptw_status_pei;
  wire core_io_ptw_status_ei;
  wire core_io_ptw_status_ps;
  wire core_io_ptw_status_s;
  wire dcache_io_cpu_req_ready;
  wire dcache_io_cpu_resp_valid;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_bits_replay;
  wire[2:0] dcache_io_cpu_resp_bits_typ;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire[63:0] dcache_io_cpu_resp_bits_data_subword;
  wire[7:0] dcache_io_cpu_resp_bits_tag;
  wire[3:0] dcache_io_cpu_resp_bits_cmd;
  wire[43:0] dcache_io_cpu_resp_bits_addr;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire dcache_io_cpu_replay_next_valid;
  wire[7:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_ptw_req_valid;
  wire[29:0] dcache_io_cpu_ptw_req_bits;
  wire dcache_io_cpu_ordered;
  wire dcache_io_mem_acquire_valid;
  wire[1:0] dcache_io_mem_acquire_bits_header_src;
  wire[1:0] dcache_io_mem_acquire_bits_header_dst;
  wire[25:0] dcache_io_mem_acquire_bits_payload_addr;
  wire[1:0] dcache_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] dcache_io_mem_acquire_bits_payload_data;
  wire[2:0] dcache_io_mem_acquire_bits_payload_a_type;
  wire[5:0] dcache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] dcache_io_mem_acquire_bits_payload_subword_addr;
  wire[3:0] dcache_io_mem_acquire_bits_payload_atomic_opcode;
  wire dcache_io_mem_grant_ready;
  wire dcache_io_mem_finish_valid;
  wire[1:0] dcache_io_mem_finish_bits_header_src;
  wire[1:0] dcache_io_mem_finish_bits_header_dst;
  wire[2:0] dcache_io_mem_finish_bits_payload_master_xact_id;
  wire dcache_io_mem_probe_ready;
  wire dcache_io_mem_release_valid;
  wire[1:0] dcache_io_mem_release_bits_header_src;
  wire[1:0] dcache_io_mem_release_bits_header_dst;
  wire[25:0] dcache_io_mem_release_bits_payload_addr;
  wire[1:0] dcache_io_mem_release_bits_payload_client_xact_id;
  wire[2:0] dcache_io_mem_release_bits_payload_master_xact_id;
  wire[511:0] dcache_io_mem_release_bits_payload_data;
  wire[2:0] dcache_io_mem_release_bits_payload_r_type;


  assign io_host_debug_stats_pcr = core_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = core_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = core_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = core_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = core_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = core_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = core_io_host_pcr_req_ready;
  assign io_tilelink_release_bits_payload_r_type = dcache_io_mem_release_bits_payload_r_type;
  assign io_tilelink_release_bits_payload_data = dcache_io_mem_release_bits_payload_data;
  assign io_tilelink_release_bits_payload_master_xact_id = dcache_io_mem_release_bits_payload_master_xact_id;
  assign io_tilelink_release_bits_payload_client_xact_id = T1;
  assign T1 = T0[1'h1:1'h0];
  assign T0 = {dcache_io_mem_release_bits_payload_client_xact_id, 1'h0};
  assign io_tilelink_release_bits_payload_addr = dcache_io_mem_release_bits_payload_addr;
  assign io_tilelink_release_bits_header_dst = dcache_io_mem_release_bits_header_dst;
  assign io_tilelink_release_bits_header_src = dcache_io_mem_release_bits_header_src;
  assign io_tilelink_release_valid = dcache_io_mem_release_valid;
  assign io_tilelink_probe_ready = dcache_io_mem_probe_ready;
  assign io_tilelink_finish_bits_payload_master_xact_id = memArb_io_out_finish_bits_payload_master_xact_id;
  assign io_tilelink_finish_bits_header_dst = memArb_io_out_finish_bits_header_dst;
  assign io_tilelink_finish_bits_header_src = memArb_io_out_finish_bits_header_src;
  assign io_tilelink_finish_valid = memArb_io_out_finish_valid;
  assign io_tilelink_grant_ready = memArb_io_out_grant_ready;
  assign io_tilelink_acquire_bits_payload_atomic_opcode = memArb_io_out_acquire_bits_payload_atomic_opcode;
  assign io_tilelink_acquire_bits_payload_subword_addr = memArb_io_out_acquire_bits_payload_subword_addr;
  assign io_tilelink_acquire_bits_payload_write_mask = memArb_io_out_acquire_bits_payload_write_mask;
  assign io_tilelink_acquire_bits_payload_a_type = memArb_io_out_acquire_bits_payload_a_type;
  assign io_tilelink_acquire_bits_payload_data = memArb_io_out_acquire_bits_payload_data;
  assign io_tilelink_acquire_bits_payload_client_xact_id = memArb_io_out_acquire_bits_payload_client_xact_id;
  assign io_tilelink_acquire_bits_payload_addr = memArb_io_out_acquire_bits_payload_addr;
  assign io_tilelink_acquire_bits_header_dst = memArb_io_out_acquire_bits_header_dst;
  assign io_tilelink_acquire_bits_header_src = memArb_io_out_acquire_bits_header_src;
  assign io_tilelink_acquire_valid = memArb_io_out_acquire_valid;
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_index( icache_io_cpu_btb_resp_bits_bht_index ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_index( core_io_imem_btb_update_bits_prediction_bits_bht_index ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_cpu_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_cpu_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_incorrectTarget( core_io_imem_btb_update_bits_incorrectTarget ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_cpu_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_0_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_0_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_0_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_0_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_0_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_0_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_0_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_0_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_0_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_0_sret ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_mem_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_1_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_1_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcArb_io_mem_req_valid ),
       .io_cpu_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_cpu_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_cpu_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_1_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_1_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_1_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_1_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_1_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_1_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_1_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_1_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_1_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_1_sret ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_mem_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_mem_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_mem_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( dcache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( dcache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( dcache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_0_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_0_finish_ready ),
       .io_mem_finish_valid( dcache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( io_tilelink_probe_valid ),
       .io_mem_probe_bits_header_src( io_tilelink_probe_bits_header_src ),
       .io_mem_probe_bits_header_dst( io_tilelink_probe_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( io_tilelink_probe_bits_payload_addr ),
       .io_mem_probe_bits_payload_master_xact_id( io_tilelink_probe_bits_payload_master_xact_id ),
       .io_mem_probe_bits_payload_p_type( io_tilelink_probe_bits_payload_p_type ),
       .io_mem_release_ready( io_tilelink_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_header_src( dcache_io_mem_release_bits_header_src ),
       .io_mem_release_bits_header_dst( dcache_io_mem_release_bits_header_dst ),
       .io_mem_release_bits_payload_addr( dcache_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( dcache_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_master_xact_id( dcache_io_mem_release_bits_payload_master_xact_id ),
       .io_mem_release_bits_payload_data( dcache_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( dcache_io_mem_release_bits_payload_r_type )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_requestor_1_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_requestor_1_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_requestor_1_status_ip( ptw_io_requestor_1_status_ip ),
       .io_requestor_1_status_im( ptw_io_requestor_1_status_im ),
       .io_requestor_1_status_zero( ptw_io_requestor_1_status_zero ),
       .io_requestor_1_status_er( ptw_io_requestor_1_status_er ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_requestor_1_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_requestor_1_status_ef( ptw_io_requestor_1_status_ef ),
       .io_requestor_1_status_pei( ptw_io_requestor_1_status_pei ),
       .io_requestor_1_status_ei( ptw_io_requestor_1_status_ei ),
       .io_requestor_1_status_ps( ptw_io_requestor_1_status_ps ),
       .io_requestor_1_status_s( ptw_io_requestor_1_status_s ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_1_sret( ptw_io_requestor_1_sret ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_requestor_0_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_requestor_0_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_requestor_0_status_ip( ptw_io_requestor_0_status_ip ),
       .io_requestor_0_status_im( ptw_io_requestor_0_status_im ),
       .io_requestor_0_status_zero( ptw_io_requestor_0_status_zero ),
       .io_requestor_0_status_er( ptw_io_requestor_0_status_er ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_requestor_0_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_requestor_0_status_ef( ptw_io_requestor_0_status_ef ),
       .io_requestor_0_status_pei( ptw_io_requestor_0_status_pei ),
       .io_requestor_0_status_ei( ptw_io_requestor_0_status_ei ),
       .io_requestor_0_status_ps( ptw_io_requestor_0_status_ps ),
       .io_requestor_0_status_s( ptw_io_requestor_0_status_s ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_requestor_0_sret( ptw_io_requestor_0_sret ),
       .io_mem_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_data(  )
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_mem_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       //.io_mem_ptw_req_valid(  )
       //.io_mem_ptw_req_bits(  )
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_sret( core_io_ptw_sret ),
       .io_dpath_status_ip( core_io_ptw_status_ip ),
       .io_dpath_status_im( core_io_ptw_status_im ),
       .io_dpath_status_zero( core_io_ptw_status_zero ),
       .io_dpath_status_er( core_io_ptw_status_er ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_s64( core_io_ptw_status_s64 ),
       .io_dpath_status_u64( core_io_ptw_status_u64 ),
       .io_dpath_status_ef( core_io_ptw_status_ef ),
       .io_dpath_status_pei( core_io_ptw_status_pei ),
       .io_dpath_status_ei( core_io_ptw_status_ei ),
       .io_dpath_status_ps( core_io_ptw_status_ps ),
       .io_dpath_status_s( core_io_ptw_status_s )
  );
  Core core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( core_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( core_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( core_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( core_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( core_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( core_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( core_io_host_debug_stats_pcr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_index( icache_io_cpu_btb_resp_bits_bht_index ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_index( core_io_imem_btb_update_bits_prediction_bits_bht_index ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_imem_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_incorrectTarget( core_io_imem_btb_update_bits_incorrectTarget ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_imem_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_dmem_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       //.io_dmem_ptw_req_valid(  )
       //.io_dmem_ptw_req_bits(  )
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( dcArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_sret( core_io_ptw_sret ),
       .io_ptw_status_ip( core_io_ptw_status_ip ),
       .io_ptw_status_im( core_io_ptw_status_im ),
       .io_ptw_status_zero( core_io_ptw_status_zero ),
       .io_ptw_status_er( core_io_ptw_status_er ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_s64( core_io_ptw_status_s64 ),
       .io_ptw_status_u64( core_io_ptw_status_u64 ),
       .io_ptw_status_ef( core_io_ptw_status_ef ),
       .io_ptw_status_pei( core_io_ptw_status_pei ),
       .io_ptw_status_ei( core_io_ptw_status_ei ),
       .io_ptw_status_ps( core_io_ptw_status_ps ),
       .io_ptw_status_s( core_io_ptw_status_s )
       //.io_rocc_cmd_ready(  )
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       //.io_rocc_resp_valid(  )
       //.io_rocc_resp_bits_rd(  )
       //.io_rocc_resp_bits_data(  )
       //.io_rocc_mem_req_ready(  )
       //.io_rocc_mem_req_valid(  )
       //.io_rocc_mem_req_bits_kill(  )
       //.io_rocc_mem_req_bits_typ(  )
       //.io_rocc_mem_req_bits_phys(  )
       //.io_rocc_mem_req_bits_addr(  )
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_req_bits_tag(  )
       //.io_rocc_mem_req_bits_cmd(  )
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_ptw_req_ready(  )
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       //.io_rocc_mem_ptw_resp_valid(  )
       //.io_rocc_mem_ptw_resp_bits_error(  )
       //.io_rocc_mem_ptw_resp_bits_ppn(  )
       //.io_rocc_mem_ptw_resp_bits_perm(  )
       //.io_rocc_mem_ptw_status_ip(  )
       //.io_rocc_mem_ptw_status_im(  )
       //.io_rocc_mem_ptw_status_zero(  )
       //.io_rocc_mem_ptw_status_er(  )
       //.io_rocc_mem_ptw_status_vm(  )
       //.io_rocc_mem_ptw_status_s64(  )
       //.io_rocc_mem_ptw_status_u64(  )
       //.io_rocc_mem_ptw_status_ef(  )
       //.io_rocc_mem_ptw_status_pei(  )
       //.io_rocc_mem_ptw_status_ei(  )
       //.io_rocc_mem_ptw_status_ps(  )
       //.io_rocc_mem_ptw_status_s(  )
       //.io_rocc_mem_ptw_invalidate(  )
       //.io_rocc_mem_ptw_sret(  )
       //.io_rocc_mem_ordered(  )
       //.io_rocc_busy(  )
       //.io_rocc_s(  )
       //.io_rocc_interrupt(  )
       //.io_rocc_imem_acquire_ready(  )
       //.io_rocc_imem_acquire_valid(  )
       //.io_rocc_imem_acquire_bits_header_src(  )
       //.io_rocc_imem_acquire_bits_header_dst(  )
       //.io_rocc_imem_acquire_bits_payload_addr(  )
       //.io_rocc_imem_acquire_bits_payload_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_payload_data(  )
       //.io_rocc_imem_acquire_bits_payload_a_type(  )
       //.io_rocc_imem_acquire_bits_payload_write_mask(  )
       //.io_rocc_imem_acquire_bits_payload_subword_addr(  )
       //.io_rocc_imem_acquire_bits_payload_atomic_opcode(  )
       //.io_rocc_imem_grant_ready(  )
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       //.io_rocc_imem_finish_valid(  )
       //.io_rocc_imem_finish_bits_header_src(  )
       //.io_rocc_imem_finish_bits_header_dst(  )
       //.io_rocc_imem_finish_bits_payload_master_xact_id(  )
       //.io_rocc_iptw_req_ready(  )
       //.io_rocc_iptw_req_valid(  )
       //.io_rocc_iptw_req_bits(  )
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       //.io_rocc_dptw_req_valid(  )
       //.io_rocc_dptw_req_bits(  )
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       //.io_rocc_pptw_req_valid(  )
       //.io_rocc_pptw_req_bits(  )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );
  `ifndef SYNTHESIS
    assign core.io_dmem_ptw_req_valid = {1{$random}};
    assign core.io_dmem_ptw_req_bits = {1{$random}};
    assign core.io_rocc_cmd_ready = {1{$random}};
    assign core.io_rocc_resp_valid = {1{$random}};
    assign core.io_rocc_resp_bits_rd = {1{$random}};
    assign core.io_rocc_resp_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_valid = {1{$random}};
    assign core.io_rocc_mem_req_bits_kill = {1{$random}};
    assign core.io_rocc_mem_req_bits_typ = {1{$random}};
    assign core.io_rocc_mem_req_bits_phys = {1{$random}};
    assign core.io_rocc_mem_req_bits_addr = {2{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_cmd = {1{$random}};
    assign core.io_rocc_mem_ptw_req_ready = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_valid = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_error = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_ppn = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_perm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ip = {1{$random}};
    assign core.io_rocc_mem_ptw_status_im = {1{$random}};
    assign core.io_rocc_mem_ptw_status_zero = {1{$random}};
    assign core.io_rocc_mem_ptw_status_er = {1{$random}};
    assign core.io_rocc_mem_ptw_status_vm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_u64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ef = {1{$random}};
    assign core.io_rocc_mem_ptw_status_pei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ps = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s = {1{$random}};
    assign core.io_rocc_mem_ptw_invalidate = {1{$random}};
    assign core.io_rocc_mem_ptw_sret = {1{$random}};
    assign core.io_rocc_busy = {1{$random}};
    assign core.io_rocc_interrupt = {1{$random}};
    assign core.io_rocc_imem_acquire_valid = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_client_xact_id = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_data = {16{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_a_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_write_mask = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_subword_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_atomic_opcode = {1{$random}};
    assign core.io_rocc_imem_grant_ready = {1{$random}};
    assign core.io_rocc_imem_finish_valid = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_finish_bits_payload_master_xact_id = {1{$random}};
    assign core.io_rocc_iptw_req_valid = {1{$random}};
    assign core.io_rocc_iptw_req_bits = {1{$random}};
    assign core.io_rocc_dptw_req_valid = {1{$random}};
    assign core.io_rocc_dptw_req_bits = {1{$random}};
    assign core.io_rocc_pptw_req_valid = {1{$random}};
    assign core.io_rocc_pptw_req_bits = {1{$random}};
  `endif
  HellaCacheArbiter dcArb(.clk(clk),
       .io_requestor_1_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_requestor_1_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_requestor_1_ptw_req_ready(  )
       //.io_requestor_1_ptw_req_valid(  )
       //.io_requestor_1_ptw_req_bits(  )
       //.io_requestor_1_ptw_resp_valid(  )
       //.io_requestor_1_ptw_resp_bits_error(  )
       //.io_requestor_1_ptw_resp_bits_ppn(  )
       //.io_requestor_1_ptw_resp_bits_perm(  )
       //.io_requestor_1_ptw_status_ip(  )
       //.io_requestor_1_ptw_status_im(  )
       //.io_requestor_1_ptw_status_zero(  )
       //.io_requestor_1_ptw_status_er(  )
       //.io_requestor_1_ptw_status_vm(  )
       //.io_requestor_1_ptw_status_s64(  )
       //.io_requestor_1_ptw_status_u64(  )
       //.io_requestor_1_ptw_status_ef(  )
       //.io_requestor_1_ptw_status_pei(  )
       //.io_requestor_1_ptw_status_ei(  )
       //.io_requestor_1_ptw_status_ps(  )
       //.io_requestor_1_ptw_status_s(  )
       //.io_requestor_1_ptw_invalidate(  )
       //.io_requestor_1_ptw_sret(  )
       .io_requestor_1_ordered( dcArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_data(  )
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_requestor_0_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_requestor_0_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_ptw_req_ready(  )
       //.io_requestor_0_ptw_req_valid(  )
       //.io_requestor_0_ptw_req_bits(  )
       //.io_requestor_0_ptw_resp_valid(  )
       //.io_requestor_0_ptw_resp_bits_error(  )
       //.io_requestor_0_ptw_resp_bits_ppn(  )
       //.io_requestor_0_ptw_resp_bits_perm(  )
       //.io_requestor_0_ptw_status_ip(  )
       //.io_requestor_0_ptw_status_im(  )
       //.io_requestor_0_ptw_status_zero(  )
       //.io_requestor_0_ptw_status_er(  )
       //.io_requestor_0_ptw_status_vm(  )
       //.io_requestor_0_ptw_status_s64(  )
       //.io_requestor_0_ptw_status_u64(  )
       //.io_requestor_0_ptw_status_ef(  )
       //.io_requestor_0_ptw_status_pei(  )
       //.io_requestor_0_ptw_status_ei(  )
       //.io_requestor_0_ptw_status_ps(  )
       //.io_requestor_0_ptw_status_s(  )
       //.io_requestor_0_ptw_invalidate(  )
       //.io_requestor_0_ptw_sret(  )
       .io_requestor_0_ordered( dcArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcArb_io_mem_req_valid ),
       .io_mem_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_mem_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       .io_mem_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_mem_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
  `ifndef SYNTHESIS
    assign dcArb.io_requestor_0_req_bits_data = {2{$random}};
    assign dcArb.io_requestor_0_req_bits_tag = {1{$random}};
  `endif
  UncachedTileLinkIOArbiterThatAppendsArbiterId memArb(.clk(clk), .reset(reset),
       .io_in_1_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_in_1_acquire_bits_header_src(  )
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_in_1_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_in_1_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_in_1_grant_ready( icache_io_mem_grant_ready ),
       .io_in_1_grant_valid( memArb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( memArb_io_in_1_finish_ready ),
       .io_in_1_finish_valid( icache_io_mem_finish_valid ),
       .io_in_1_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_in_1_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_in_1_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_in_0_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_in_0_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_in_0_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_write_mask( dcache_io_mem_acquire_bits_payload_write_mask ),
       .io_in_0_acquire_bits_payload_subword_addr( dcache_io_mem_acquire_bits_payload_subword_addr ),
       .io_in_0_acquire_bits_payload_atomic_opcode( dcache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_in_0_grant_ready( dcache_io_mem_grant_ready ),
       .io_in_0_grant_valid( memArb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( memArb_io_in_0_finish_ready ),
       .io_in_0_finish_valid( dcache_io_mem_finish_valid ),
       .io_in_0_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_in_0_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_in_0_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_acquire_ready( io_tilelink_acquire_ready ),
       .io_out_acquire_valid( memArb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( memArb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( memArb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( memArb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( memArb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( memArb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_a_type( memArb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_write_mask( memArb_io_out_acquire_bits_payload_write_mask ),
       .io_out_acquire_bits_payload_subword_addr( memArb_io_out_acquire_bits_payload_subword_addr ),
       .io_out_acquire_bits_payload_atomic_opcode( memArb_io_out_acquire_bits_payload_atomic_opcode ),
       .io_out_grant_ready( memArb_io_out_grant_ready ),
       .io_out_grant_valid( io_tilelink_grant_valid ),
       .io_out_grant_bits_header_src( io_tilelink_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_tilelink_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_tilelink_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_tilelink_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_tilelink_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_g_type( io_tilelink_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_tilelink_finish_ready ),
       .io_out_finish_valid( memArb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( memArb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( memArb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( memArb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign memArb.io_in_1_acquire_bits_header_src = {1{$random}};
    assign memArb.io_in_1_acquire_bits_header_dst = {1{$random}};
  `endif
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [1:0] io_enq_bits_client_xact_id,
    input [511:0] io_enq_bits_data,
    input [2:0] io_enq_bits_a_type,
    input [5:0] io_enq_bits_write_mask,
    input [2:0] io_enq_bits_subword_addr,
    input [3:0] io_enq_bits_atomic_opcode,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[1:0] io_deq_bits_client_xact_id,
    output[511:0] io_deq_bits_data,
    output[2:0] io_deq_bits_a_type,
    output[5:0] io_deq_bits_write_mask,
    output[2:0] io_deq_bits_subword_addr,
    output[3:0] io_deq_bits_atomic_opcode,
    output io_count
);

  wire T21;
  wire[1:0] T0;
  reg  full;
  wire T22;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[3:0] T3;
  wire[555:0] T4;
  reg [555:0] ram [0:0];
  wire[555:0] T5;
  wire[555:0] T6;
  wire[555:0] T7;
  wire[15:0] T8;
  wire[6:0] T9;
  wire[8:0] T10;
  wire[539:0] T11;
  wire[513:0] T12;
  wire[2:0] T13;
  wire[5:0] T14;
  wire[2:0] T15;
  wire[511:0] T16;
  wire[1:0] T17;
  wire[25:0] T18;
  wire T19;
  wire empty;
  wire T20;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {18{$random}};
  end
`endif

  assign io_count = T21;
  assign T21 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T22 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_atomic_opcode = T3;
  assign T3 = T4[2'h3:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = {io_enq_bits_subword_addr, io_enq_bits_atomic_opcode};
  assign T10 = {io_enq_bits_a_type, io_enq_bits_write_mask};
  assign T11 = {io_enq_bits_addr, T12};
  assign T12 = {io_enq_bits_client_xact_id, io_enq_bits_data};
  assign io_deq_bits_subword_addr = T13;
  assign T13 = T4[3'h6:3'h4];
  assign io_deq_bits_write_mask = T14;
  assign T14 = T4[4'hc:3'h7];
  assign io_deq_bits_a_type = T15;
  assign T15 = T4[4'hf:4'hd];
  assign io_deq_bits_data = T16;
  assign T16 = T4[10'h20f:5'h10];
  assign io_deq_bits_client_xact_id = T17;
  assign T17 = T4[10'h211:10'h210];
  assign io_deq_bits_addr = T18;
  assign T18 = T4[10'h22b:10'h212];
  assign io_deq_valid = T19;
  assign T19 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module HTIF(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    output io_cpu_0_reset,
    //output io_cpu_0_id
    input  io_cpu_0_pcr_req_ready,
    output io_cpu_0_pcr_req_valid,
    output io_cpu_0_pcr_req_bits_rw,
    output[4:0] io_cpu_0_pcr_req_bits_addr,
    output[63:0] io_cpu_0_pcr_req_bits_data,
    output io_cpu_0_pcr_rep_ready,
    input  io_cpu_0_pcr_rep_valid,
    input [63:0] io_cpu_0_pcr_rep_bits,
    output io_cpu_0_ipi_req_ready,
    input  io_cpu_0_ipi_req_valid,
    input  io_cpu_0_ipi_req_bits,
    input  io_cpu_0_ipi_rep_ready,
    output io_cpu_0_ipi_rep_valid,
    //output io_cpu_0_ipi_rep_bits
    input  io_cpu_0_debug_stats_pcr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    //output[1:0] io_mem_finish_bits_header_src
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [2:0] io_mem_probe_bits_payload_master_xact_id,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    //output[1:0] io_mem_release_bits_header_src
    //output[1:0] io_mem_release_bits_header_dst
    output[25:0] io_mem_release_bits_payload_addr,
    output[1:0] io_mem_release_bits_payload_client_xact_id,
    output[2:0] io_mem_release_bits_payload_master_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    //input [63:0] io_scr_rdata_1
    //input [63:0] io_scr_rdata_0
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire[3:0] T347;
  wire[3:0] T348;
  wire[3:0] T349;
  wire T350;
  reg [3:0] cmd;
  wire[3:0] T20;
  wire[3:0] next_cmd;
  wire[63:0] rx_shifter_in;
  wire[47:0] T30;
  reg [63:0] rx_shifter;
  wire[63:0] T31;
  wire T59;
  wire T21;
  wire T22;
  reg [14:0] rx_count;
  wire[14:0] T337;
  wire[14:0] T23;
  wire[14:0] T24;
  wire[14:0] T25;
  wire T26;
  wire T27;
  wire[12:0] T338;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T28;
  wire[11:0] T29;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire nack;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire bad_mem_packet;
  wire T44;
  wire[2:0] T45;
  reg [39:0] addr;
  wire[39:0] T46;
  wire[39:0] T47;
  wire[39:0] T48;
  wire[39:0] T49;
  wire T96;
  wire T97;
  reg [3:0] state;
  wire[3:0] T336;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  wire[3:0] rx_cmd;
  wire T60;
  wire[12:0] rx_word_count;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire rx_done;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire T69;
  wire[12:0] T340;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire rx_word_done;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  reg  mem_acked;
  wire T341;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire[3:0] T88;
  wire T89;
  wire T90;
  reg [8:0] pos;
  wire[8:0] T91;
  wire[8:0] T92;
  wire[8:0] T93;
  wire[8:0] T94;
  wire T95;
  wire[3:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T112;
  wire T113;
  wire T114;
  wire[4:0] pcr_addr;
  wire T115;
  wire T116;
  wire[1:0] pcr_coreid;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[12:0] tx_word_count;
  reg [14:0] tx_count;
  wire[14:0] T339;
  wire[14:0] T55;
  wire[14:0] T56;
  wire[14:0] T57;
  wire T58;
  wire T102;
  wire tx_done;
  wire T103;
  wire T104;
  wire T105;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T106;
  wire T107;
  wire T108;
  wire[12:0] T342;
  wire T109;
  wire T110;
  wire[1:0] tx_subword_count;
  wire T111;
  wire[2:0] T351;
  wire[2:0] T352;
  wire[2:0] T353;
  wire[5:0] T354;
  wire[5:0] T355;
  wire[5:0] T356;
  wire[2:0] T357;
  wire[2:0] T358;
  wire[2:0] T359;
  wire[511:0] T360;
  wire[511:0] T361;
  wire[511:0] T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[25:0] T366;
  wire[25:0] T367;
  wire[25:0] T368;
  wire[36:0] init_addr;
  wire[39:0] T369;
  wire[25:0] T370;
  wire[25:0] T371;
  wire T372;
  wire T373;
  wire T374;
  wire[63:0] pcr_wdata;
  reg [63:0] packet_ram [7:0];
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire T3;
  wire[63:0] T121;
  wire[63:0] T122;
  wire T123;
  wire T124;
  wire[63:0] T125;
  wire[63:0] T126;
  wire T127;
  wire T128;
  wire[63:0] T129;
  wire[63:0] T130;
  wire T131;
  wire T132;
  wire[63:0] T133;
  wire[63:0] T134;
  wire T135;
  wire T136;
  wire[63:0] T137;
  wire[63:0] T138;
  wire T139;
  wire T140;
  wire[63:0] T141;
  wire[63:0] T142;
  wire T143;
  wire T144;
  wire[63:0] T145;
  wire[63:0] T146;
  wire T147;
  wire T148;
  wire[63:0] T149;
  wire T150;
  wire[2:0] T151;
  wire[2:0] T152;
  wire[5:0] T153;
  wire[5:0] scr_addr;
  wire T154;
  wire T155;
  reg [2:0] mem_gxid;
  wire[2:0] T156;
  reg [1:0] mem_gsrc;
  wire[1:0] T157;
  wire T158;
  reg  mem_needs_ack;
  wire T159;
  wire T160;
  wire T161;
  wire[511:0] mem_req_data;
  wire[447:0] T162;
  wire[383:0] T163;
  wire[319:0] T164;
  wire[255:0] T165;
  wire[191:0] T166;
  wire[127:0] T167;
  wire[63:0] T168;
  wire[63:0] T169;
  wire[63:0] T170;
  wire[63:0] T171;
  wire[63:0] T172;
  wire[63:0] T173;
  wire[63:0] T174;
  wire[63:0] T175;
  reg  R176;
  wire T343;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  reg  R186;
  wire T344;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire[15:0] T345;
  wire[63:0] T191;
  wire[5:0] T192;
  wire[1:0] T193;
  wire[63:0] tx_data;
  wire[63:0] T194;
  wire[63:0] T195;
  reg [63:0] pcrReadData;
  wire[63:0] T196;
  wire[63:0] T197;
  wire[63:0] T198;
  wire[63:0] T346;
  wire[63:0] T199;
  wire[63:0] T200;
  wire[63:0] T201;
  wire[63:0] T202;
  wire[63:0] T203;
  wire[63:0] T204;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T205;
  wire[5:0] T206;
  wire[63:0] T207;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T208;
  wire T209;
  wire[63:0] T210;
  wire[63:0] T211;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T212;
  wire[63:0] T213;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T214;
  wire T215;
  wire T216;
  wire[63:0] T217;
  wire[63:0] T218;
  wire[63:0] T219;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T220;
  wire[63:0] T221;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T222;
  wire T223;
  wire[63:0] T224;
  wire[63:0] T225;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T226;
  wire[63:0] T227;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire[63:0] T232;
  wire[63:0] T233;
  wire[63:0] T234;
  wire[63:0] T235;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T236;
  wire[63:0] T237;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T238;
  wire T239;
  wire[63:0] T240;
  wire[63:0] T241;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T242;
  wire[63:0] T243;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T244;
  wire T245;
  wire T246;
  wire[63:0] T247;
  wire[63:0] T248;
  wire[63:0] T249;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T250;
  wire[63:0] T251;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T252;
  wire T253;
  wire[63:0] T254;
  wire[63:0] T255;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T256;
  wire[63:0] T257;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire[63:0] T263;
  wire[63:0] T264;
  wire[63:0] T265;
  wire[63:0] T266;
  wire[63:0] T267;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T268;
  wire[63:0] T269;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T270;
  wire T271;
  wire[63:0] T272;
  wire[63:0] T273;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T274;
  wire[63:0] T275;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T276;
  wire T277;
  wire T278;
  wire[63:0] T279;
  wire[63:0] T280;
  wire[63:0] T281;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T282;
  wire[63:0] T283;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T284;
  wire T285;
  wire[63:0] T286;
  wire[63:0] T287;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T288;
  wire[63:0] T289;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire[63:0] T294;
  wire[63:0] T295;
  wire[63:0] T296;
  wire[63:0] T297;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T298;
  wire[63:0] T299;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T300;
  wire T301;
  wire[63:0] T302;
  wire[63:0] T303;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T304;
  wire[63:0] T305;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T306;
  wire T307;
  wire T308;
  wire[63:0] T309;
  wire[63:0] T310;
  wire[63:0] T311;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T312;
  wire[63:0] T313;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T314;
  wire T315;
  wire[63:0] T316;
  wire[63:0] T317;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T318;
  wire[63:0] T319;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[63:0] tx_header;
  wire[15:0] T329;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T330;
  reg [7:0] seqno;
  wire[7:0] T331;
  wire[7:0] T332;
  wire T333;
  wire T334;
  wire T335;
  wire acq_q_io_enq_ready;
  wire acq_q_io_deq_valid;
  wire[25:0] acq_q_io_deq_bits_addr;
  wire[1:0] acq_q_io_deq_bits_client_xact_id;
  wire[2:0] acq_q_io_deq_bits_a_type;
  wire[5:0] acq_q_io_deq_bits_write_mask;
  wire[2:0] acq_q_io_deq_bits_subword_addr;
  wire[3:0] acq_q_io_deq_bits_atomic_opcode;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cmd = {1{$random}};
    rx_shifter = {2{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    addr = {2{$random}};
    state = {1{$random}};
    mem_acked = {1{$random}};
    pos = {1{$random}};
    tx_count = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    mem_gxid = {1{$random}};
    mem_gsrc = {1{$random}};
    mem_needs_ack = {1{$random}};
    R176 = {1{$random}};
    R186 = {1{$random}};
    pcrReadData = {2{$random}};
    seqno = {1{$random}};
  end
`endif

  assign T347 = T350 ? T349 : T348;
  assign T348 = 4'h0;
  assign T349 = 4'h0;
  assign T350 = cmd == 4'h1;
  assign T20 = T21 ? next_cmd : cmd;
  assign next_cmd = rx_shifter_in[2'h3:1'h0];
  assign rx_shifter_in = {io_host_in_bits, T30};
  assign T30 = rx_shifter[6'h3f:5'h10];
  assign T31 = T59 ? rx_shifter_in : rx_shifter;
  assign T59 = io_host_in_valid & io_host_in_ready;
  assign T21 = T59 & T22;
  assign T22 = rx_count == 15'h3;
  assign T337 = reset ? 15'h0 : T23;
  assign T23 = T26 ? 15'h0 : T24;
  assign T24 = T59 ? T25 : rx_count;
  assign T25 = rx_count + 15'h1;
  assign T26 = T102 & T27;
  assign T27 = tx_word_count == T338;
  assign T338 = {1'h0, tx_size};
  assign tx_size = T32 ? size : 12'h0;
  assign T28 = T21 ? T29 : size;
  assign T29 = rx_shifter_in[4'hf:3'h4];
  assign T32 = T38 & T33;
  assign T33 = T35 | T34;
  assign T34 = cmd == 4'h3;
  assign T35 = T37 | T36;
  assign T36 = cmd == 4'h2;
  assign T37 = cmd == 4'h0;
  assign T38 = nack ^ 1'h1;
  assign nack = T52 ? bad_mem_packet : T39;
  assign T39 = T41 ? T40 : 1'h1;
  assign T40 = size != 12'h1;
  assign T41 = T43 | T42;
  assign T42 = cmd == 4'h3;
  assign T43 = cmd == 4'h2;
  assign bad_mem_packet = T50 | T44;
  assign T44 = T45 != 3'h0;
  assign T45 = addr[2'h2:1'h0];
  assign T46 = T96 ? T49 : T47;
  assign T47 = T21 ? T48 : addr;
  assign T48 = rx_shifter_in[6'h3f:5'h18];
  assign T49 = addr + 40'h8;
  assign T96 = T97 & io_mem_finish_ready;
  assign T97 = state == 4'h7;
  assign T336 = reset ? 4'h0 : T4;
  assign T4 = T118 ? 4'h8 : T5;
  assign T5 = io_cpu_0_pcr_rep_valid ? 4'h8 : T6;
  assign T6 = T113 ? 4'h8 : T7;
  assign T7 = T112 ? 4'h2 : T8;
  assign T8 = T102 ? T98 : T9;
  assign T9 = T96 ? T88 : T10;
  assign T10 = T87 ? 4'h7 : T11;
  assign T11 = T81 ? 4'h7 : T12;
  assign T12 = T79 ? 4'h5 : T13;
  assign T13 = T77 ? 4'h6 : T14;
  assign T14 = T64 ? T15 : state;
  assign T15 = T63 ? 4'h3 : T16;
  assign T16 = T62 ? 4'h4 : T17;
  assign T17 = T18 ? 4'h1 : 4'h8;
  assign T18 = T61 | T19;
  assign T19 = rx_cmd == 4'h3;
  assign rx_cmd = T60 ? next_cmd : cmd;
  assign T60 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T61 = rx_cmd == 4'h2;
  assign T62 = rx_cmd == 4'h1;
  assign T63 = rx_cmd == 4'h0;
  assign T64 = T76 & rx_done;
  assign rx_done = rx_word_done & T65;
  assign T65 = T73 ? T70 : T66;
  assign T66 = T69 | T67;
  assign T67 = T68 == 3'h0;
  assign T68 = rx_word_count[2'h2:1'h0];
  assign T69 = rx_word_count == T340;
  assign T340 = {1'h0, size};
  assign T70 = T72 & T71;
  assign T71 = next_cmd != 4'h3;
  assign T72 = next_cmd != 4'h1;
  assign T73 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T74;
  assign T74 = T75 == 2'h3;
  assign T75 = rx_count[1'h1:1'h0];
  assign T76 = state == 4'h0;
  assign T77 = T78 & acq_q_io_enq_ready;
  assign T78 = state == 4'h4;
  assign T79 = T80 & acq_q_io_enq_ready;
  assign T80 = state == 4'h3;
  assign T81 = T86 & mem_acked;
  assign T341 = reset ? 1'h0 : T82;
  assign T82 = T85 ? 1'h0 : T83;
  assign T83 = T81 ? 1'h0 : T84;
  assign T84 = io_mem_grant_valid ? 1'h1 : mem_acked;
  assign T85 = state == 4'h5;
  assign T86 = state == 4'h6;
  assign T87 = T85 & io_mem_grant_valid;
  assign T88 = T89 ? 4'h8 : 4'h0;
  assign T89 = T95 | T90;
  assign T90 = pos == 9'h1;
  assign T91 = T96 ? T94 : T92;
  assign T92 = T21 ? T93 : pos;
  assign T93 = rx_shifter_in[4'hf:3'h7];
  assign T94 = pos - 9'h1;
  assign T95 = cmd == 4'h0;
  assign T98 = T99 ? 4'h3 : 4'h0;
  assign T99 = T101 & T100;
  assign T100 = pos != 9'h0;
  assign T101 = cmd == 4'h0;
  assign T112 = io_cpu_0_pcr_req_valid & io_cpu_0_pcr_req_ready;
  assign T113 = T115 & T114;
  assign T114 = pcr_addr == 5'h1d;
  assign pcr_addr = addr[3'h4:1'h0];
  assign T115 = T117 & T116;
  assign T116 = pcr_coreid == 2'h0;
  assign pcr_coreid = addr[5'h15:5'h14];
  assign T117 = state == 4'h1;
  assign T118 = T120 & T119;
  assign T119 = pcr_coreid == 2'h3;
  assign T120 = state == 4'h1;
  assign T50 = T51 != 3'h0;
  assign T51 = size[2'h2:1'h0];
  assign T52 = T54 | T53;
  assign T53 = cmd == 4'h1;
  assign T54 = cmd == 4'h0;
  assign tx_word_count = tx_count[4'he:2'h2];
  assign T339 = reset ? 15'h0 : T55;
  assign T55 = T26 ? 15'h0 : T56;
  assign T56 = T58 ? T57 : tx_count;
  assign T57 = tx_count + 15'h1;
  assign T58 = io_host_out_valid & io_host_out_ready;
  assign T102 = T111 & tx_done;
  assign tx_done = T109 & T103;
  assign T103 = T108 | T104;
  assign T104 = T107 & T105;
  assign T105 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T106 - 3'h1;
  assign T106 = tx_word_count[2'h2:1'h0];
  assign T107 = 13'h0 < tx_word_count;
  assign T108 = tx_word_count == T342;
  assign T342 = {1'h0, tx_size};
  assign T109 = io_host_out_ready & T110;
  assign T110 = tx_subword_count == 2'h3;
  assign tx_subword_count = tx_count[1'h1:1'h0];
  assign T111 = state == 4'h8;
  assign T351 = T350 ? T353 : T352;
  assign T352 = 3'h0;
  assign T353 = 3'h0;
  assign T354 = T350 ? T356 : T355;
  assign T355 = 6'h0;
  assign T356 = 6'h0;
  assign T357 = T350 ? T359 : T358;
  assign T358 = 3'h2;
  assign T359 = 3'h3;
  assign T360 = T350 ? T362 : T361;
  assign T361 = 512'h0;
  assign T362 = 512'h0;
  assign T363 = T350 ? T365 : T364;
  assign T364 = 2'h0;
  assign T365 = 2'h0;
  assign T366 = T350 ? T370 : T367;
  assign T367 = T368;
  assign T368 = init_addr[5'h19:1'h0];
  assign init_addr = T369 >> 2'h3;
  assign T369 = addr;
  assign T370 = T371;
  assign T371 = init_addr[5'h19:1'h0];
  assign T372 = T374 | T373;
  assign T373 = state == 4'h4;
  assign T374 = state == 4'h3;
  assign io_scr_wdata = pcr_wdata;
  assign pcr_wdata = packet_ram[3'h0];
  assign T1 = io_mem_grant_bits_payload_data[9'h1ff:9'h1c0];
  assign T2 = T3 & io_mem_grant_valid;
  assign T3 = state == 4'h5;
  assign T122 = io_mem_grant_bits_payload_data[9'h1bf:9'h180];
  assign T123 = T124 & io_mem_grant_valid;
  assign T124 = state == 4'h5;
  assign T126 = io_mem_grant_bits_payload_data[9'h17f:9'h140];
  assign T127 = T128 & io_mem_grant_valid;
  assign T128 = state == 4'h5;
  assign T130 = io_mem_grant_bits_payload_data[9'h13f:9'h100];
  assign T131 = T132 & io_mem_grant_valid;
  assign T132 = state == 4'h5;
  assign T134 = io_mem_grant_bits_payload_data[8'hff:8'hc0];
  assign T135 = T136 & io_mem_grant_valid;
  assign T136 = state == 4'h5;
  assign T138 = io_mem_grant_bits_payload_data[8'hbf:8'h80];
  assign T139 = T140 & io_mem_grant_valid;
  assign T140 = state == 4'h5;
  assign T142 = io_mem_grant_bits_payload_data[7'h7f:7'h40];
  assign T143 = T144 & io_mem_grant_valid;
  assign T144 = state == 4'h5;
  assign T146 = io_mem_grant_bits_payload_data[6'h3f:1'h0];
  assign T147 = T148 & io_mem_grant_valid;
  assign T148 = state == 4'h5;
  assign T150 = rx_word_done & io_host_in_ready;
  assign T151 = T152 - 3'h1;
  assign T152 = rx_word_count[2'h2:1'h0];
  assign io_scr_waddr = T153;
  assign T153 = scr_addr;
  assign scr_addr = addr[3'h5:1'h0];
  assign io_scr_wen = T154;
  assign T154 = T118 ? T155 : 1'h0;
  assign T155 = cmd == 4'h3;
  assign io_mem_release_valid = 1'h0;
  assign io_mem_probe_ready = 1'h0;
  assign io_mem_finish_bits_payload_master_xact_id = mem_gxid;
  assign T156 = io_mem_grant_valid ? io_mem_grant_bits_payload_master_xact_id : mem_gxid;
  assign io_mem_finish_bits_header_dst = mem_gsrc;
  assign T157 = io_mem_grant_valid ? io_mem_grant_bits_header_src : mem_gsrc;
  assign io_mem_finish_valid = T158;
  assign T158 = T161 & mem_needs_ack;
  assign T159 = io_mem_grant_valid ? T160 : mem_needs_ack;
  assign T160 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T161 = state == 4'h7;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_payload_atomic_opcode = acq_q_io_deq_bits_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = acq_q_io_deq_bits_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = acq_q_io_deq_bits_write_mask;
  assign io_mem_acquire_bits_payload_a_type = acq_q_io_deq_bits_a_type;
  assign io_mem_acquire_bits_payload_data = mem_req_data;
  assign mem_req_data = {T175, T162};
  assign T162 = {T174, T163};
  assign T163 = {T173, T164};
  assign T164 = {T172, T165};
  assign T165 = {T171, T166};
  assign T166 = {T170, T167};
  assign T167 = {T169, T168};
  assign T168 = packet_ram[3'h0];
  assign T169 = packet_ram[3'h1];
  assign T170 = packet_ram[3'h2];
  assign T171 = packet_ram[3'h3];
  assign T172 = packet_ram[3'h4];
  assign T173 = packet_ram[3'h5];
  assign T174 = packet_ram[3'h6];
  assign T175 = packet_ram[3'h7];
  assign io_mem_acquire_bits_payload_client_xact_id = acq_q_io_deq_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = acq_q_io_deq_bits_addr;
  assign io_mem_acquire_bits_header_dst = 2'h0;
  assign io_mem_acquire_bits_header_src = 2'h2;
  assign io_mem_acquire_valid = acq_q_io_deq_valid;
  assign io_cpu_0_ipi_rep_valid = R176;
  assign T343 = reset ? 1'h0 : T177;
  assign T177 = T179 ? 1'h1 : T178;
  assign T178 = io_cpu_0_ipi_rep_ready ? 1'h0 : R176;
  assign T179 = io_cpu_0_ipi_req_valid & T180;
  assign T180 = io_cpu_0_ipi_req_bits == 1'h0;
  assign io_cpu_0_ipi_req_ready = 1'h1;
  assign io_cpu_0_pcr_rep_ready = 1'h1;
  assign io_cpu_0_pcr_req_bits_data = pcr_wdata;
  assign io_cpu_0_pcr_req_bits_addr = pcr_addr;
  assign io_cpu_0_pcr_req_bits_rw = T181;
  assign T181 = cmd == 4'h3;
  assign io_cpu_0_pcr_req_valid = T182;
  assign T182 = T184 & T183;
  assign T183 = pcr_addr != 5'h1d;
  assign T184 = T185 & T116;
  assign T185 = state == 4'h1;
  assign io_cpu_0_reset = R186;
  assign T344 = reset ? 1'h1 : T187;
  assign T187 = T189 ? T188 : R186;
  assign T188 = pcr_wdata[1'h0:1'h0];
  assign T189 = T113 & T190;
  assign T190 = cmd == 4'h3;
  assign io_host_debug_stats_pcr = io_cpu_0_debug_stats_pcr;
  assign io_host_out_bits = T345;
  assign T345 = T191[4'hf:1'h0];
  assign T191 = tx_data >> T192;
  assign T192 = {T193, 4'h0};
  assign T193 = tx_count[1'h1:1'h0];
  assign tx_data = T333 ? tx_header : T194;
  assign T194 = T326 ? pcrReadData : T195;
  assign T195 = packet_ram[packet_ram_raddr];
  assign T196 = T118 ? T199 : T197;
  assign T197 = io_cpu_0_pcr_rep_valid ? io_cpu_0_pcr_rep_bits : T198;
  assign T198 = T113 ? T346 : pcrReadData;
  assign T346 = {63'h0, R186};
  assign T199 = T325 ? T263 : T200;
  assign T200 = T262 ? T232 : T201;
  assign T201 = T231 ? T217 : T202;
  assign T202 = T216 ? T210 : T203;
  assign T203 = T209 ? T207 : T204;
  assign T204 = T205 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = 64'h1;
  assign scr_rdata_1 = 64'h1000;
  assign T205 = T206[1'h0:1'h0];
  assign T206 = scr_addr;
  assign T207 = T208 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T208 = T206[1'h0:1'h0];
  assign T209 = T206[1'h1:1'h1];
  assign T210 = T215 ? T213 : T211;
  assign T211 = T212 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T212 = T206[1'h0:1'h0];
  assign T213 = T214 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T214 = T206[1'h0:1'h0];
  assign T215 = T206[1'h1:1'h1];
  assign T216 = T206[2'h2:2'h2];
  assign T217 = T230 ? T224 : T218;
  assign T218 = T223 ? T221 : T219;
  assign T219 = T220 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T220 = T206[1'h0:1'h0];
  assign T221 = T222 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T222 = T206[1'h0:1'h0];
  assign T223 = T206[1'h1:1'h1];
  assign T224 = T229 ? T227 : T225;
  assign T225 = T226 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T226 = T206[1'h0:1'h0];
  assign T227 = T228 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T228 = T206[1'h0:1'h0];
  assign T229 = T206[1'h1:1'h1];
  assign T230 = T206[2'h2:2'h2];
  assign T231 = T206[2'h3:2'h3];
  assign T232 = T261 ? T247 : T233;
  assign T233 = T246 ? T240 : T234;
  assign T234 = T239 ? T237 : T235;
  assign T235 = T236 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T236 = T206[1'h0:1'h0];
  assign T237 = T238 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T238 = T206[1'h0:1'h0];
  assign T239 = T206[1'h1:1'h1];
  assign T240 = T245 ? T243 : T241;
  assign T241 = T242 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T242 = T206[1'h0:1'h0];
  assign T243 = T244 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T244 = T206[1'h0:1'h0];
  assign T245 = T206[1'h1:1'h1];
  assign T246 = T206[2'h2:2'h2];
  assign T247 = T260 ? T254 : T248;
  assign T248 = T253 ? T251 : T249;
  assign T249 = T250 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T250 = T206[1'h0:1'h0];
  assign T251 = T252 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T252 = T206[1'h0:1'h0];
  assign T253 = T206[1'h1:1'h1];
  assign T254 = T259 ? T257 : T255;
  assign T255 = T256 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T256 = T206[1'h0:1'h0];
  assign T257 = T258 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T258 = T206[1'h0:1'h0];
  assign T259 = T206[1'h1:1'h1];
  assign T260 = T206[2'h2:2'h2];
  assign T261 = T206[2'h3:2'h3];
  assign T262 = T206[3'h4:3'h4];
  assign T263 = T324 ? T294 : T264;
  assign T264 = T293 ? T279 : T265;
  assign T265 = T278 ? T272 : T266;
  assign T266 = T271 ? T269 : T267;
  assign T267 = T268 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T268 = T206[1'h0:1'h0];
  assign T269 = T270 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T270 = T206[1'h0:1'h0];
  assign T271 = T206[1'h1:1'h1];
  assign T272 = T277 ? T275 : T273;
  assign T273 = T274 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T274 = T206[1'h0:1'h0];
  assign T275 = T276 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T276 = T206[1'h0:1'h0];
  assign T277 = T206[1'h1:1'h1];
  assign T278 = T206[2'h2:2'h2];
  assign T279 = T292 ? T286 : T280;
  assign T280 = T285 ? T283 : T281;
  assign T281 = T282 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T282 = T206[1'h0:1'h0];
  assign T283 = T284 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T284 = T206[1'h0:1'h0];
  assign T285 = T206[1'h1:1'h1];
  assign T286 = T291 ? T289 : T287;
  assign T287 = T288 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T288 = T206[1'h0:1'h0];
  assign T289 = T290 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T290 = T206[1'h0:1'h0];
  assign T291 = T206[1'h1:1'h1];
  assign T292 = T206[2'h2:2'h2];
  assign T293 = T206[2'h3:2'h3];
  assign T294 = T323 ? T309 : T295;
  assign T295 = T308 ? T302 : T296;
  assign T296 = T301 ? T299 : T297;
  assign T297 = T298 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T298 = T206[1'h0:1'h0];
  assign T299 = T300 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T300 = T206[1'h0:1'h0];
  assign T301 = T206[1'h1:1'h1];
  assign T302 = T307 ? T305 : T303;
  assign T303 = T304 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T304 = T206[1'h0:1'h0];
  assign T305 = T306 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T306 = T206[1'h0:1'h0];
  assign T307 = T206[1'h1:1'h1];
  assign T308 = T206[2'h2:2'h2];
  assign T309 = T322 ? T316 : T310;
  assign T310 = T315 ? T313 : T311;
  assign T311 = T312 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T312 = T206[1'h0:1'h0];
  assign T313 = T314 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T314 = T206[1'h0:1'h0];
  assign T315 = T206[1'h1:1'h1];
  assign T316 = T321 ? T319 : T317;
  assign T317 = T318 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T318 = T206[1'h0:1'h0];
  assign T319 = T320 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T320 = T206[1'h0:1'h0];
  assign T321 = T206[1'h1:1'h1];
  assign T322 = T206[2'h2:2'h2];
  assign T323 = T206[2'h3:2'h3];
  assign T324 = T206[3'h4:3'h4];
  assign T325 = T206[3'h5:3'h5];
  assign T326 = T328 | T327;
  assign T327 = cmd == 4'h3;
  assign T328 = cmd == 4'h2;
  assign tx_header = {T330, T329};
  assign T329 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T330 = {addr, seqno};
  assign T331 = T21 ? T332 : seqno;
  assign T332 = rx_shifter_in[5'h17:5'h10];
  assign T333 = tx_word_count == 13'h0;
  assign io_host_out_valid = T334;
  assign T334 = state == 4'h8;
  assign io_host_in_ready = T335;
  assign T335 = state == 4'h0;
  Queue_8 acq_q(.clk(clk), .reset(reset),
       .io_enq_ready( acq_q_io_enq_ready ),
       .io_enq_valid( T372 ),
       .io_enq_bits_addr( T366 ),
       .io_enq_bits_client_xact_id( T363 ),
       .io_enq_bits_data( T360 ),
       .io_enq_bits_a_type( T357 ),
       .io_enq_bits_write_mask( T354 ),
       .io_enq_bits_subword_addr( T351 ),
       .io_enq_bits_atomic_opcode( T347 ),
       .io_deq_ready( io_mem_acquire_ready ),
       .io_deq_valid( acq_q_io_deq_valid ),
       .io_deq_bits_addr( acq_q_io_deq_bits_addr ),
       .io_deq_bits_client_xact_id( acq_q_io_deq_bits_client_xact_id ),
       //.io_deq_bits_data(  )
       .io_deq_bits_a_type( acq_q_io_deq_bits_a_type ),
       .io_deq_bits_write_mask( acq_q_io_deq_bits_write_mask ),
       .io_deq_bits_subword_addr( acq_q_io_deq_bits_subword_addr ),
       .io_deq_bits_atomic_opcode( acq_q_io_deq_bits_atomic_opcode )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T21) begin
      cmd <= next_cmd;
    end
    if(T59) begin
      rx_shifter <= rx_shifter_in;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T26) begin
      rx_count <= 15'h0;
    end else if(T59) begin
      rx_count <= T25;
    end
    if(T21) begin
      size <= T29;
    end
    if(T96) begin
      addr <= T49;
    end else if(T21) begin
      addr <= T48;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T118) begin
      state <= 4'h8;
    end else if(io_cpu_0_pcr_rep_valid) begin
      state <= 4'h8;
    end else if(T113) begin
      state <= 4'h8;
    end else if(T112) begin
      state <= 4'h2;
    end else if(T102) begin
      state <= T98;
    end else if(T96) begin
      state <= T88;
    end else if(T87) begin
      state <= 4'h7;
    end else if(T81) begin
      state <= 4'h7;
    end else if(T79) begin
      state <= 4'h5;
    end else if(T77) begin
      state <= 4'h6;
    end else if(T64) begin
      state <= T15;
    end
    if(reset) begin
      mem_acked <= 1'h0;
    end else if(T85) begin
      mem_acked <= 1'h0;
    end else if(T81) begin
      mem_acked <= 1'h0;
    end else if(io_mem_grant_valid) begin
      mem_acked <= 1'h1;
    end
    if(T96) begin
      pos <= T94;
    end else if(T21) begin
      pos <= T93;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T26) begin
      tx_count <= 15'h0;
    end else if(T58) begin
      tx_count <= T57;
    end
    if (T2)
      packet_ram[3'h7] <= T1;
    if (T123)
      packet_ram[3'h6] <= T122;
    if (T127)
      packet_ram[3'h5] <= T126;
    if (T131)
      packet_ram[3'h4] <= T130;
    if (T135)
      packet_ram[3'h3] <= T134;
    if (T139)
      packet_ram[3'h2] <= T138;
    if (T143)
      packet_ram[3'h1] <= T142;
    if (T147)
      packet_ram[3'h0] <= T146;
    if (T150)
      packet_ram[T151] <= rx_shifter_in;
    if(io_mem_grant_valid) begin
      mem_gxid <= io_mem_grant_bits_payload_master_xact_id;
    end
    if(io_mem_grant_valid) begin
      mem_gsrc <= io_mem_grant_bits_header_src;
    end
    if(io_mem_grant_valid) begin
      mem_needs_ack <= T160;
    end
    if(reset) begin
      R176 <= 1'h0;
    end else if(T179) begin
      R176 <= 1'h1;
    end else if(io_cpu_0_ipi_rep_ready) begin
      R176 <= 1'h0;
    end
    if(reset) begin
      R186 <= 1'h1;
    end else if(T189) begin
      R186 <= T188;
    end
    if(T118) begin
      pcrReadData <= T199;
    end else if(io_cpu_0_pcr_rep_valid) begin
      pcrReadData <= io_cpu_0_pcr_rep_bits;
    end else if(T113) begin
      pcrReadData <= T346;
    end
    if(T21) begin
      seqno <= T332;
    end
  end
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T83;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire[5:0] T19;
  wire[5:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire T25;
  wire T26;
  wire[511:0] T27;
  wire[511:0] T28;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire[25:0] T35;
  wire[25:0] T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T83 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_atomic_opcode = T10;
  assign T10 = T14 ? io_in_2_bits_payload_atomic_opcode : T11;
  assign T11 = T12 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_subword_addr = T15;
  assign T15 = T18 ? io_in_2_bits_payload_subword_addr : T16;
  assign T16 = T17 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_write_mask = T19;
  assign T19 = T22 ? io_in_2_bits_payload_write_mask : T20;
  assign T20 = T21 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T23;
  assign T23 = T26 ? io_in_2_bits_payload_a_type : T24;
  assign T24 = T25 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_payload_data = T27;
  assign T27 = T30 ? io_in_2_bits_payload_data : T28;
  assign T28 = T29 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T31;
  assign T31 = T34 ? io_in_2_bits_payload_client_xact_id : T32;
  assign T32 = T33 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_out_bits_payload_addr = T35;
  assign T35 = T38 ? io_in_2_bits_payload_addr : T36;
  assign T36 = T37 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T37 = T13[1'h0:1'h0];
  assign T38 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T39;
  assign T39 = T42 ? io_in_2_bits_header_dst : T40;
  assign T40 = T41 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T41 = T13[1'h0:1'h0];
  assign T42 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T43;
  assign T43 = T46 ? io_in_2_bits_header_src : T44;
  assign T44 = T45 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T45 = T13[1'h0:1'h0];
  assign T46 = T13[1'h1:1'h1];
  assign io_out_valid = T47;
  assign T47 = T50 ? io_in_2_valid : T48;
  assign T48 = T49 ? io_in_1_valid : io_in_0_valid;
  assign T49 = T13[1'h0:1'h0];
  assign T50 = T13[1'h1:1'h1];
  assign io_in_0_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T62 | T53;
  assign T53 = T54 ^ 1'h1;
  assign T54 = T57 | T55;
  assign T55 = io_in_2_valid & T56;
  assign T56 = last_grant < 2'h2;
  assign T57 = T60 | T58;
  assign T58 = io_in_1_valid & T59;
  assign T59 = last_grant < 2'h1;
  assign T60 = io_in_0_valid & T61;
  assign T61 = last_grant < 2'h0;
  assign T62 = last_grant < 2'h0;
  assign io_in_1_ready = T63;
  assign T63 = T64 & io_out_ready;
  assign T64 = T69 | T65;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_0_valid;
  assign T67 = T68 | T55;
  assign T68 = T60 | T58;
  assign T69 = T71 & T70;
  assign T70 = last_grant < 2'h1;
  assign T71 = T60 ^ 1'h1;
  assign io_in_2_ready = T72;
  assign T72 = T73 & io_out_ready;
  assign T73 = T79 | T74;
  assign T74 = T75 ^ 1'h1;
  assign T75 = T76 | io_in_1_valid;
  assign T76 = T77 | io_in_0_valid;
  assign T77 = T78 | T55;
  assign T78 = T60 | T58;
  assign T79 = T81 & T80;
  assign T80 = last_grant < 2'h2;
  assign T81 = T82 ^ 1'h1;
  assign T82 = T60 | T58;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_a_type,
    output[5:0] io_out_2_bits_payload_write_mask,
    output[2:0] io_out_2_bits_payload_subword_addr,
    output[3:0] io_out_2_bits_payload_atomic_opcode,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_a_type,
    output[5:0] io_out_1_bits_payload_write_mask,
    output[2:0] io_out_1_bits_payload_subword_addr,
    output[3:0] io_out_1_bits_payload_atomic_opcode,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_a_type,
    output[5:0] io_out_0_bits_payload_write_mask,
    output[2:0] io_out_0_bits_payload_subword_addr,
    output[3:0] io_out_0_bits_payload_atomic_opcode
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_0_io_in_2_ready;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire LockingRRArbiter_0_io_out_valid;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_a_type;
  wire[5:0] LockingRRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_subword_addr;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_a_type;
  wire[5:0] LockingRRArbiter_1_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_subword_addr;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_atomic_opcode;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire LockingRRArbiter_2_io_out_valid;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_a_type;
  wire[5:0] LockingRRArbiter_2_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_subword_addr;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_atomic_opcode;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_atomic_opcode = LockingRRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_0_bits_payload_subword_addr = LockingRRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_0_bits_payload_write_mask = LockingRRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_0_bits_payload_a_type = LockingRRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_atomic_opcode = LockingRRArbiter_1_io_out_bits_payload_atomic_opcode;
  assign io_out_1_bits_payload_subword_addr = LockingRRArbiter_1_io_out_bits_payload_subword_addr;
  assign io_out_1_bits_payload_write_mask = LockingRRArbiter_1_io_out_bits_payload_write_mask;
  assign io_out_1_bits_payload_a_type = LockingRRArbiter_1_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_atomic_opcode = LockingRRArbiter_2_io_out_bits_payload_atomic_opcode;
  assign io_out_2_bits_payload_subword_addr = LockingRRArbiter_2_io_out_bits_payload_subword_addr;
  assign io_out_2_bits_payload_write_mask = LockingRRArbiter_2_io_out_bits_payload_write_mask;
  assign io_out_2_bits_payload_a_type = LockingRRArbiter_2_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_2_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_2_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_1_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_0_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_2_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_1_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_0_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_2_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_1_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_0_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_0 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_1_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_1_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_1_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_1_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_2_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_2_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_2_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_2_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_r_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T75;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[511:0] T15;
  wire[511:0] T16;
  wire T17;
  wire T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire[25:0] T27;
  wire[25:0] T28;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T75 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_r_type = T10;
  assign T10 = T14 ? io_in_2_bits_payload_r_type : T11;
  assign T11 = T12 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_data = T15;
  assign T15 = T18 ? io_in_2_bits_payload_data : T16;
  assign T16 = T17 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T19;
  assign T19 = T22 ? io_in_2_bits_payload_master_xact_id : T20;
  assign T20 = T21 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T23;
  assign T23 = T26 ? io_in_2_bits_payload_client_xact_id : T24;
  assign T24 = T25 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_payload_addr = T27;
  assign T27 = T30 ? io_in_2_bits_payload_addr : T28;
  assign T28 = T29 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T31;
  assign T31 = T34 ? io_in_2_bits_header_dst : T32;
  assign T32 = T33 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T35;
  assign T35 = T38 ? io_in_2_bits_header_src : T36;
  assign T36 = T37 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T37 = T13[1'h0:1'h0];
  assign T38 = T13[1'h1:1'h1];
  assign io_out_valid = T39;
  assign T39 = T42 ? io_in_2_valid : T40;
  assign T40 = T41 ? io_in_1_valid : io_in_0_valid;
  assign T41 = T13[1'h0:1'h0];
  assign T42 = T13[1'h1:1'h1];
  assign io_in_0_ready = T43;
  assign T43 = T44 & io_out_ready;
  assign T44 = T54 | T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T49 | T47;
  assign T47 = io_in_2_valid & T48;
  assign T48 = last_grant < 2'h2;
  assign T49 = T52 | T50;
  assign T50 = io_in_1_valid & T51;
  assign T51 = last_grant < 2'h1;
  assign T52 = io_in_0_valid & T53;
  assign T53 = last_grant < 2'h0;
  assign T54 = last_grant < 2'h0;
  assign io_in_1_ready = T55;
  assign T55 = T56 & io_out_ready;
  assign T56 = T61 | T57;
  assign T57 = T58 ^ 1'h1;
  assign T58 = T59 | io_in_0_valid;
  assign T59 = T60 | T47;
  assign T60 = T52 | T50;
  assign T61 = T63 & T62;
  assign T62 = last_grant < 2'h1;
  assign T63 = T52 ^ 1'h1;
  assign io_in_2_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T71 | T66;
  assign T66 = T67 ^ 1'h1;
  assign T67 = T68 | io_in_1_valid;
  assign T68 = T69 | io_in_0_valid;
  assign T69 = T70 | T47;
  assign T70 = T52 | T50;
  assign T71 = T73 & T72;
  assign T72 = last_grant < 2'h2;
  assign T73 = T74 ^ 1'h1;
  assign T74 = T52 | T50;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_r_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_r_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_r_type
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_3_io_in_2_ready;
  wire LockingRRArbiter_3_io_in_1_ready;
  wire LockingRRArbiter_3_io_in_0_ready;
  wire LockingRRArbiter_3_io_out_valid;
  wire[1:0] LockingRRArbiter_3_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_3_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_3_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_3_io_out_bits_payload_master_xact_id;
  wire[511:0] LockingRRArbiter_3_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_3_io_out_bits_payload_r_type;
  wire LockingRRArbiter_4_io_in_2_ready;
  wire LockingRRArbiter_4_io_in_1_ready;
  wire LockingRRArbiter_4_io_in_0_ready;
  wire LockingRRArbiter_4_io_out_valid;
  wire[1:0] LockingRRArbiter_4_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_4_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_4_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_4_io_out_bits_payload_master_xact_id;
  wire[511:0] LockingRRArbiter_4_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_4_io_out_bits_payload_r_type;
  wire LockingRRArbiter_5_io_in_2_ready;
  wire LockingRRArbiter_5_io_in_1_ready;
  wire LockingRRArbiter_5_io_in_0_ready;
  wire LockingRRArbiter_5_io_out_valid;
  wire[1:0] LockingRRArbiter_5_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_5_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_5_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_5_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_5_io_out_bits_payload_master_xact_id;
  wire[511:0] LockingRRArbiter_5_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_5_io_out_bits_payload_r_type;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_r_type = LockingRRArbiter_3_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_3_io_out_bits_payload_data;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_3_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_3_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_3_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_3_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_3_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_3_io_out_valid;
  assign io_out_1_bits_payload_r_type = LockingRRArbiter_4_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_4_io_out_bits_payload_data;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_4_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_4_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_4_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_4_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_4_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_4_io_out_valid;
  assign io_out_2_bits_payload_r_type = LockingRRArbiter_5_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_5_io_out_bits_payload_data;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_5_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_5_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_5_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_5_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_5_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_5_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_5_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_4_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_3_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_5_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_4_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_3_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_5_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_4_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_3_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_1 LockingRRArbiter_3(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_3_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_3_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_3_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_3_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_3_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_4(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_4_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_4_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_4_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_4_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_4_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_4_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_4_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_4_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_4_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_4_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_4_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_5(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_5_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_5_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_5_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_5_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_5_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_5_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_5_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_5_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_5_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_5_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_5_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_out_bits_payload_p_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T67;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire[25:0] T19;
  wire[25:0] T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T67 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_p_type = T10;
  assign T10 = T14 ? io_in_2_bits_payload_p_type : T11;
  assign T11 = T12 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T15;
  assign T15 = T18 ? io_in_2_bits_payload_master_xact_id : T16;
  assign T16 = T17 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_addr = T19;
  assign T19 = T22 ? io_in_2_bits_payload_addr : T20;
  assign T20 = T21 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T23;
  assign T23 = T26 ? io_in_2_bits_header_dst : T24;
  assign T24 = T25 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T27;
  assign T27 = T30 ? io_in_2_bits_header_src : T28;
  assign T28 = T29 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_valid = T31;
  assign T31 = T34 ? io_in_2_valid : T32;
  assign T32 = T33 ? io_in_1_valid : io_in_0_valid;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_in_0_ready = T35;
  assign T35 = T36 & io_out_ready;
  assign T36 = T46 | T37;
  assign T37 = T38 ^ 1'h1;
  assign T38 = T41 | T39;
  assign T39 = io_in_2_valid & T40;
  assign T40 = last_grant < 2'h2;
  assign T41 = T44 | T42;
  assign T42 = io_in_1_valid & T43;
  assign T43 = last_grant < 2'h1;
  assign T44 = io_in_0_valid & T45;
  assign T45 = last_grant < 2'h0;
  assign T46 = last_grant < 2'h0;
  assign io_in_1_ready = T47;
  assign T47 = T48 & io_out_ready;
  assign T48 = T53 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_0_valid;
  assign T51 = T52 | T39;
  assign T52 = T44 | T42;
  assign T53 = T55 & T54;
  assign T54 = last_grant < 2'h1;
  assign T55 = T44 ^ 1'h1;
  assign io_in_2_ready = T56;
  assign T56 = T57 & io_out_ready;
  assign T57 = T63 | T58;
  assign T58 = T59 ^ 1'h1;
  assign T59 = T60 | io_in_1_valid;
  assign T60 = T61 | io_in_0_valid;
  assign T61 = T62 | T39;
  assign T62 = T44 | T42;
  assign T63 = T65 & T64;
  assign T64 = last_grant < 2'h2;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T44 | T42;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output[1:0] io_out_2_bits_payload_p_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output[1:0] io_out_1_bits_payload_p_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output[1:0] io_out_0_bits_payload_p_type
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_6_io_in_2_ready;
  wire LockingRRArbiter_6_io_in_1_ready;
  wire LockingRRArbiter_6_io_in_0_ready;
  wire LockingRRArbiter_6_io_out_valid;
  wire[1:0] LockingRRArbiter_6_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_6_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_6_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_6_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_6_io_out_bits_payload_p_type;
  wire LockingRRArbiter_7_io_in_2_ready;
  wire LockingRRArbiter_7_io_in_1_ready;
  wire LockingRRArbiter_7_io_in_0_ready;
  wire LockingRRArbiter_7_io_out_valid;
  wire[1:0] LockingRRArbiter_7_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_7_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_7_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_7_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_7_io_out_bits_payload_p_type;
  wire LockingRRArbiter_8_io_in_2_ready;
  wire LockingRRArbiter_8_io_in_1_ready;
  wire LockingRRArbiter_8_io_in_0_ready;
  wire LockingRRArbiter_8_io_out_valid;
  wire[1:0] LockingRRArbiter_8_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_8_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_8_io_out_bits_payload_addr;
  wire[2:0] LockingRRArbiter_8_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_8_io_out_bits_payload_p_type;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_p_type = LockingRRArbiter_6_io_out_bits_payload_p_type;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_6_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_6_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_6_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_6_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_6_io_out_valid;
  assign io_out_1_bits_payload_p_type = LockingRRArbiter_7_io_out_bits_payload_p_type;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_7_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_7_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_7_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_7_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_7_io_out_valid;
  assign io_out_2_bits_payload_p_type = LockingRRArbiter_8_io_out_bits_payload_p_type;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_8_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_8_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_8_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_8_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_8_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_8_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_7_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_6_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_8_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_7_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_6_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_8_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_7_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_6_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_2 LockingRRArbiter_6(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_6_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_6_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_6_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_6_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_6_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_6_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_6_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_6_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_6_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_7(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_7_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_7_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_7_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_7_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_7_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_7_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_7_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_7_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_7_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_8(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_8_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_8_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_8_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_8_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_8_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_8_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_8_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_8_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_8_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T71;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[511:0] T23;
  wire[511:0] T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T71 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_g_type = T10;
  assign T10 = T14 ? io_in_2_bits_payload_g_type : T11;
  assign T11 = T12 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T15;
  assign T15 = T18 ? io_in_2_bits_payload_master_xact_id : T16;
  assign T16 = T17 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T19;
  assign T19 = T22 ? io_in_2_bits_payload_client_xact_id : T20;
  assign T20 = T21 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_bits_payload_data = T23;
  assign T23 = T26 ? io_in_2_bits_payload_data : T24;
  assign T24 = T25 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T27;
  assign T27 = T30 ? io_in_2_bits_header_dst : T28;
  assign T28 = T29 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T29 = T13[1'h0:1'h0];
  assign T30 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T31;
  assign T31 = T34 ? io_in_2_bits_header_src : T32;
  assign T32 = T33 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T33 = T13[1'h0:1'h0];
  assign T34 = T13[1'h1:1'h1];
  assign io_out_valid = T35;
  assign T35 = T38 ? io_in_2_valid : T36;
  assign T36 = T37 ? io_in_1_valid : io_in_0_valid;
  assign T37 = T13[1'h0:1'h0];
  assign T38 = T13[1'h1:1'h1];
  assign io_in_0_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T50 | T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T45 | T43;
  assign T43 = io_in_2_valid & T44;
  assign T44 = last_grant < 2'h2;
  assign T45 = T48 | T46;
  assign T46 = io_in_1_valid & T47;
  assign T47 = last_grant < 2'h1;
  assign T48 = io_in_0_valid & T49;
  assign T49 = last_grant < 2'h0;
  assign T50 = last_grant < 2'h0;
  assign io_in_1_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T57 | T53;
  assign T53 = T54 ^ 1'h1;
  assign T54 = T55 | io_in_0_valid;
  assign T55 = T56 | T43;
  assign T56 = T48 | T46;
  assign T57 = T59 & T58;
  assign T58 = last_grant < 2'h1;
  assign T59 = T48 ^ 1'h1;
  assign io_in_2_ready = T60;
  assign T60 = T61 & io_out_ready;
  assign T61 = T67 | T62;
  assign T62 = T63 ^ 1'h1;
  assign T63 = T64 | io_in_1_valid;
  assign T64 = T65 | io_in_0_valid;
  assign T65 = T66 | T43;
  assign T66 = T48 | T46;
  assign T67 = T69 & T68;
  assign T68 = last_grant < 2'h2;
  assign T69 = T70 ^ 1'h1;
  assign T70 = T48 | T46;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[511:0] io_out_2_bits_payload_data,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output[3:0] io_out_2_bits_payload_g_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[511:0] io_out_1_bits_payload_data,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output[3:0] io_out_1_bits_payload_g_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[511:0] io_out_0_bits_payload_data,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output[3:0] io_out_0_bits_payload_g_type
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_9_io_in_2_ready;
  wire LockingRRArbiter_9_io_in_1_ready;
  wire LockingRRArbiter_9_io_in_0_ready;
  wire LockingRRArbiter_9_io_out_valid;
  wire[1:0] LockingRRArbiter_9_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_9_io_out_bits_header_dst;
  wire[511:0] LockingRRArbiter_9_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_9_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_9_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_9_io_out_bits_payload_g_type;
  wire LockingRRArbiter_10_io_in_2_ready;
  wire LockingRRArbiter_10_io_in_1_ready;
  wire LockingRRArbiter_10_io_in_0_ready;
  wire LockingRRArbiter_10_io_out_valid;
  wire[1:0] LockingRRArbiter_10_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_10_io_out_bits_header_dst;
  wire[511:0] LockingRRArbiter_10_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_10_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_10_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_10_io_out_bits_payload_g_type;
  wire LockingRRArbiter_11_io_in_2_ready;
  wire LockingRRArbiter_11_io_in_1_ready;
  wire LockingRRArbiter_11_io_in_0_ready;
  wire LockingRRArbiter_11_io_out_valid;
  wire[1:0] LockingRRArbiter_11_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_11_io_out_bits_header_dst;
  wire[511:0] LockingRRArbiter_11_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_11_io_out_bits_payload_client_xact_id;
  wire[2:0] LockingRRArbiter_11_io_out_bits_payload_master_xact_id;
  wire[3:0] LockingRRArbiter_11_io_out_bits_payload_g_type;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_g_type = LockingRRArbiter_9_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_9_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_9_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_data = LockingRRArbiter_9_io_out_bits_payload_data;
  assign io_out_0_bits_header_dst = LockingRRArbiter_9_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_9_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_9_io_out_valid;
  assign io_out_1_bits_payload_g_type = LockingRRArbiter_10_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_10_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_10_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_data = LockingRRArbiter_10_io_out_bits_payload_data;
  assign io_out_1_bits_header_dst = LockingRRArbiter_10_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_10_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_10_io_out_valid;
  assign io_out_2_bits_payload_g_type = LockingRRArbiter_11_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_11_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_11_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_data = LockingRRArbiter_11_io_out_bits_payload_data;
  assign io_out_2_bits_header_dst = LockingRRArbiter_11_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_11_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_11_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_11_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_10_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_9_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_11_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_10_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_9_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_11_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_10_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_9_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_3 LockingRRArbiter_9(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_9_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_9_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_9_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_9_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_9_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_9_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_9_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_9_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_9_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_9_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_10(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_10_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_10_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_10_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_10_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_10_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_10_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_10_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_10_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_10_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_10_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_11(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_11_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_11_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_11_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_11_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_11_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_11_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_11_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_11_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_11_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_11_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T59;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire[1:0] T13;
  wire T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T59 = reset ? 2'h0 : T6;
  assign T6 = T7 ? T0 : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign io_out_bits_payload_master_xact_id = T10;
  assign T10 = T14 ? io_in_2_bits_payload_master_xact_id : T11;
  assign T11 = T12 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = T0;
  assign T14 = T13[1'h1:1'h1];
  assign io_out_bits_header_dst = T15;
  assign T15 = T18 ? io_in_2_bits_header_dst : T16;
  assign T16 = T17 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T17 = T13[1'h0:1'h0];
  assign T18 = T13[1'h1:1'h1];
  assign io_out_bits_header_src = T19;
  assign T19 = T22 ? io_in_2_bits_header_src : T20;
  assign T20 = T21 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T21 = T13[1'h0:1'h0];
  assign T22 = T13[1'h1:1'h1];
  assign io_out_valid = T23;
  assign T23 = T26 ? io_in_2_valid : T24;
  assign T24 = T25 ? io_in_1_valid : io_in_0_valid;
  assign T25 = T13[1'h0:1'h0];
  assign T26 = T13[1'h1:1'h1];
  assign io_in_0_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T38 | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T33 | T31;
  assign T31 = io_in_2_valid & T32;
  assign T32 = last_grant < 2'h2;
  assign T33 = T36 | T34;
  assign T34 = io_in_1_valid & T35;
  assign T35 = last_grant < 2'h1;
  assign T36 = io_in_0_valid & T37;
  assign T37 = last_grant < 2'h0;
  assign T38 = last_grant < 2'h0;
  assign io_in_1_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T45 | T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T43 | io_in_0_valid;
  assign T43 = T44 | T31;
  assign T44 = T36 | T34;
  assign T45 = T47 & T46;
  assign T46 = last_grant < 2'h1;
  assign T47 = T36 ^ 1'h1;
  assign io_in_2_ready = T48;
  assign T48 = T49 & io_out_ready;
  assign T49 = T55 | T50;
  assign T50 = T51 ^ 1'h1;
  assign T51 = T52 | io_in_1_valid;
  assign T52 = T53 | io_in_0_valid;
  assign T53 = T54 | T31;
  assign T54 = T36 | T34;
  assign T55 = T57 & T56;
  assign T56 = last_grant < 2'h2;
  assign T57 = T58 ^ 1'h1;
  assign T58 = T36 | T34;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[2:0] io_out_0_bits_payload_master_xact_id
);

  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_12_io_in_2_ready;
  wire LockingRRArbiter_12_io_in_1_ready;
  wire LockingRRArbiter_12_io_in_0_ready;
  wire LockingRRArbiter_12_io_out_valid;
  wire[1:0] LockingRRArbiter_12_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_12_io_out_bits_header_dst;
  wire[2:0] LockingRRArbiter_12_io_out_bits_payload_master_xact_id;
  wire LockingRRArbiter_13_io_in_2_ready;
  wire LockingRRArbiter_13_io_in_1_ready;
  wire LockingRRArbiter_13_io_in_0_ready;
  wire LockingRRArbiter_13_io_out_valid;
  wire[1:0] LockingRRArbiter_13_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_13_io_out_bits_header_dst;
  wire[2:0] LockingRRArbiter_13_io_out_bits_payload_master_xact_id;
  wire LockingRRArbiter_14_io_in_2_ready;
  wire LockingRRArbiter_14_io_in_1_ready;
  wire LockingRRArbiter_14_io_in_0_ready;
  wire LockingRRArbiter_14_io_out_valid;
  wire[1:0] LockingRRArbiter_14_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_14_io_out_bits_header_dst;
  wire[2:0] LockingRRArbiter_14_io_out_bits_payload_master_xact_id;


  assign T33 = io_in_0_valid & T34;
  assign T34 = io_in_0_bits_header_dst == 2'h2;
  assign T35 = io_in_1_valid & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h2;
  assign T37 = io_in_2_valid & T38;
  assign T38 = io_in_2_bits_header_dst == 2'h2;
  assign T39 = io_in_0_valid & T40;
  assign T40 = io_in_0_bits_header_dst == 2'h1;
  assign T41 = io_in_1_valid & T42;
  assign T42 = io_in_1_bits_header_dst == 2'h1;
  assign T43 = io_in_2_valid & T44;
  assign T44 = io_in_2_bits_header_dst == 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = io_in_0_bits_header_dst == 2'h0;
  assign T47 = io_in_1_valid & T48;
  assign T48 = io_in_1_bits_header_dst == 2'h0;
  assign T49 = io_in_2_valid & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_12_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_header_dst = LockingRRArbiter_12_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_12_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_12_io_out_valid;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_13_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_header_dst = LockingRRArbiter_13_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_13_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_13_io_out_valid;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_14_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_header_dst = LockingRRArbiter_14_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_14_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_14_io_out_valid;
  assign io_in_0_ready = T0;
  assign T0 = T4 | T1;
  assign T1 = T2;
  assign T2 = LockingRRArbiter_14_io_in_0_ready & T3;
  assign T3 = io_in_0_bits_header_dst == 2'h2;
  assign T4 = T8 | T5;
  assign T5 = T6;
  assign T6 = LockingRRArbiter_13_io_in_0_ready & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = T9;
  assign T9 = LockingRRArbiter_12_io_in_0_ready & T10;
  assign T10 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T11;
  assign T11 = T15 | T12;
  assign T12 = T13;
  assign T13 = LockingRRArbiter_14_io_in_1_ready & T14;
  assign T14 = io_in_1_bits_header_dst == 2'h2;
  assign T15 = T19 | T16;
  assign T16 = T17;
  assign T17 = LockingRRArbiter_13_io_in_1_ready & T18;
  assign T18 = io_in_1_bits_header_dst == 2'h1;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_12_io_in_1_ready & T21;
  assign T21 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T22;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_14_io_in_2_ready & T25;
  assign T25 = io_in_2_bits_header_dst == 2'h2;
  assign T26 = T30 | T27;
  assign T27 = T28;
  assign T28 = LockingRRArbiter_13_io_in_2_ready & T29;
  assign T29 = io_in_2_bits_header_dst == 2'h1;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_12_io_in_2_ready & T32;
  assign T32 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_4 LockingRRArbiter_12(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_12_io_in_2_ready ),
       .io_in_2_valid( T49 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_12_io_in_1_ready ),
       .io_in_1_valid( T47 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_12_io_in_0_ready ),
       .io_in_0_valid( T45 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_12_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_12_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_12_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_12_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_13(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_13_io_in_2_ready ),
       .io_in_2_valid( T43 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_13_io_in_1_ready ),
       .io_in_1_valid( T41 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_13_io_in_0_ready ),
       .io_in_0_valid( T39 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_13_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_13_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_13_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_13_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_14(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_14_io_in_2_ready ),
       .io_in_2_valid( T37 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_14_io_in_1_ready ),
       .io_in_1_valid( T35 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_14_io_in_0_ready ),
       .io_in_0_valid( T33 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_14_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_14_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_14_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_14_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module RocketChipCrossbarNetwork(input clk, input reset,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [1:0] io_clients_1_acquire_bits_header_src,
    input [1:0] io_clients_1_acquire_bits_header_dst,
    input [25:0] io_clients_1_acquire_bits_payload_addr,
    input [1:0] io_clients_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_1_acquire_bits_payload_data,
    input [2:0] io_clients_1_acquire_bits_payload_a_type,
    input [5:0] io_clients_1_acquire_bits_payload_write_mask,
    input [2:0] io_clients_1_acquire_bits_payload_subword_addr,
    input [3:0] io_clients_1_acquire_bits_payload_atomic_opcode,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_header_src,
    output[1:0] io_clients_1_grant_bits_header_dst,
    output[511:0] io_clients_1_grant_bits_payload_data,
    output[1:0] io_clients_1_grant_bits_payload_client_xact_id,
    output[2:0] io_clients_1_grant_bits_payload_master_xact_id,
    output[3:0] io_clients_1_grant_bits_payload_g_type,
    output io_clients_1_finish_ready,
    input  io_clients_1_finish_valid,
    input [1:0] io_clients_1_finish_bits_header_src,
    input [1:0] io_clients_1_finish_bits_header_dst,
    input [2:0] io_clients_1_finish_bits_payload_master_xact_id,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[1:0] io_clients_1_probe_bits_header_src,
    output[1:0] io_clients_1_probe_bits_header_dst,
    output[25:0] io_clients_1_probe_bits_payload_addr,
    output[2:0] io_clients_1_probe_bits_payload_master_xact_id,
    output[1:0] io_clients_1_probe_bits_payload_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [1:0] io_clients_1_release_bits_header_src,
    input [1:0] io_clients_1_release_bits_header_dst,
    input [25:0] io_clients_1_release_bits_payload_addr,
    input [1:0] io_clients_1_release_bits_payload_client_xact_id,
    input [2:0] io_clients_1_release_bits_payload_master_xact_id,
    input [511:0] io_clients_1_release_bits_payload_data,
    input [2:0] io_clients_1_release_bits_payload_r_type,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [1:0] io_clients_0_acquire_bits_header_src,
    input [1:0] io_clients_0_acquire_bits_header_dst,
    input [25:0] io_clients_0_acquire_bits_payload_addr,
    input [1:0] io_clients_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_0_acquire_bits_payload_data,
    input [2:0] io_clients_0_acquire_bits_payload_a_type,
    input [5:0] io_clients_0_acquire_bits_payload_write_mask,
    input [2:0] io_clients_0_acquire_bits_payload_subword_addr,
    input [3:0] io_clients_0_acquire_bits_payload_atomic_opcode,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_header_src,
    output[1:0] io_clients_0_grant_bits_header_dst,
    output[511:0] io_clients_0_grant_bits_payload_data,
    output[1:0] io_clients_0_grant_bits_payload_client_xact_id,
    output[2:0] io_clients_0_grant_bits_payload_master_xact_id,
    output[3:0] io_clients_0_grant_bits_payload_g_type,
    output io_clients_0_finish_ready,
    input  io_clients_0_finish_valid,
    input [1:0] io_clients_0_finish_bits_header_src,
    input [1:0] io_clients_0_finish_bits_header_dst,
    input [2:0] io_clients_0_finish_bits_payload_master_xact_id,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[1:0] io_clients_0_probe_bits_header_src,
    output[1:0] io_clients_0_probe_bits_header_dst,
    output[25:0] io_clients_0_probe_bits_payload_addr,
    output[2:0] io_clients_0_probe_bits_payload_master_xact_id,
    output[1:0] io_clients_0_probe_bits_payload_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [1:0] io_clients_0_release_bits_header_src,
    input [1:0] io_clients_0_release_bits_header_dst,
    input [25:0] io_clients_0_release_bits_payload_addr,
    input [1:0] io_clients_0_release_bits_payload_client_xact_id,
    input [2:0] io_clients_0_release_bits_payload_master_xact_id,
    input [511:0] io_clients_0_release_bits_payload_data,
    input [2:0] io_clients_0_release_bits_payload_r_type,
    input  io_masters_0_acquire_ready,
    output io_masters_0_acquire_valid,
    output[1:0] io_masters_0_acquire_bits_header_src,
    output[1:0] io_masters_0_acquire_bits_header_dst,
    output[25:0] io_masters_0_acquire_bits_payload_addr,
    output[1:0] io_masters_0_acquire_bits_payload_client_xact_id,
    output[511:0] io_masters_0_acquire_bits_payload_data,
    output[2:0] io_masters_0_acquire_bits_payload_a_type,
    output[5:0] io_masters_0_acquire_bits_payload_write_mask,
    output[2:0] io_masters_0_acquire_bits_payload_subword_addr,
    output[3:0] io_masters_0_acquire_bits_payload_atomic_opcode,
    output io_masters_0_grant_ready,
    input  io_masters_0_grant_valid,
    input [1:0] io_masters_0_grant_bits_header_src,
    input [1:0] io_masters_0_grant_bits_header_dst,
    input [511:0] io_masters_0_grant_bits_payload_data,
    input [1:0] io_masters_0_grant_bits_payload_client_xact_id,
    input [2:0] io_masters_0_grant_bits_payload_master_xact_id,
    input [3:0] io_masters_0_grant_bits_payload_g_type,
    input  io_masters_0_finish_ready,
    output io_masters_0_finish_valid,
    output[1:0] io_masters_0_finish_bits_header_src,
    output[1:0] io_masters_0_finish_bits_header_dst,
    output[2:0] io_masters_0_finish_bits_payload_master_xact_id,
    output io_masters_0_probe_ready,
    input  io_masters_0_probe_valid,
    input [1:0] io_masters_0_probe_bits_header_src,
    input [1:0] io_masters_0_probe_bits_header_dst,
    input [25:0] io_masters_0_probe_bits_payload_addr,
    input [2:0] io_masters_0_probe_bits_payload_master_xact_id,
    input [1:0] io_masters_0_probe_bits_payload_p_type,
    input  io_masters_0_release_ready,
    output io_masters_0_release_valid,
    output[1:0] io_masters_0_release_bits_header_src,
    output[1:0] io_masters_0_release_bits_header_dst,
    output[25:0] io_masters_0_release_bits_payload_addr,
    output[1:0] io_masters_0_release_bits_payload_client_xact_id,
    output[2:0] io_masters_0_release_bits_payload_master_xact_id,
    output[511:0] io_masters_0_release_bits_payload_data,
    output[2:0] io_masters_0_release_bits_payload_r_type
);

  wire T63;
  wire[2:0] T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[2:0] T69;
  wire[1:0] T70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[3:0] T76;
  wire[2:0] T77;
  wire[1:0] T78;
  wire[511:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[2:0] T87;
  wire[25:0] T88;
  wire[1:0] T89;
  wire[1:0] T90;
  wire[1:0] T91;
  wire T92;
  wire T93;
  wire[2:0] T94;
  wire[511:0] T95;
  wire[2:0] T96;
  wire[1:0] T97;
  wire[25:0] T98;
  wire[1:0] T99;
  wire[1:0] T100;
  wire[1:0] T101;
  wire T102;
  wire[2:0] T103;
  wire[511:0] T104;
  wire[2:0] T105;
  wire[1:0] T106;
  wire[25:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire[1:0] T110;
  wire T111;
  wire T112;
  wire[3:0] T113;
  wire[2:0] T114;
  wire[5:0] T115;
  wire[2:0] T116;
  wire[511:0] T117;
  wire[1:0] T118;
  wire[25:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire T123;
  wire[3:0] T124;
  wire[2:0] T125;
  wire[5:0] T126;
  wire[2:0] T127;
  wire[511:0] T128;
  wire[1:0] T129;
  wire[25:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire T134;
  wire[2:0] T0;
  wire[511:0] T1;
  wire[2:0] T2;
  wire[1:0] T3;
  wire[25:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire[3:0] T16;
  wire[2:0] T17;
  wire[5:0] T18;
  wire[2:0] T19;
  wire[511:0] T20;
  wire[1:0] T21;
  wire[25:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire[2:0] T29;
  wire[25:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire[3:0] T36;
  wire[2:0] T37;
  wire[1:0] T38;
  wire[511:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[1:0] T46;
  wire[2:0] T47;
  wire[25:0] T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[3:0] T54;
  wire[2:0] T55;
  wire[1:0] T56;
  wire[511:0] T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire acqNet_io_in_2_ready;
  wire acqNet_io_in_1_ready;
  wire acqNet_io_out_0_valid;
  wire[1:0] acqNet_io_out_0_bits_header_src;
  wire[1:0] acqNet_io_out_0_bits_header_dst;
  wire[25:0] acqNet_io_out_0_bits_payload_addr;
  wire[1:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire[511:0] acqNet_io_out_0_bits_payload_data;
  wire[2:0] acqNet_io_out_0_bits_payload_a_type;
  wire[5:0] acqNet_io_out_0_bits_payload_write_mask;
  wire[2:0] acqNet_io_out_0_bits_payload_subword_addr;
  wire[3:0] acqNet_io_out_0_bits_payload_atomic_opcode;
  wire relNet_io_in_2_ready;
  wire relNet_io_in_1_ready;
  wire relNet_io_out_0_valid;
  wire[1:0] relNet_io_out_0_bits_header_src;
  wire[1:0] relNet_io_out_0_bits_header_dst;
  wire[25:0] relNet_io_out_0_bits_payload_addr;
  wire[1:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire[2:0] relNet_io_out_0_bits_payload_master_xact_id;
  wire[511:0] relNet_io_out_0_bits_payload_data;
  wire[2:0] relNet_io_out_0_bits_payload_r_type;
  wire prbNet_io_in_0_ready;
  wire prbNet_io_out_2_valid;
  wire[1:0] prbNet_io_out_2_bits_header_src;
  wire[1:0] prbNet_io_out_2_bits_header_dst;
  wire[25:0] prbNet_io_out_2_bits_payload_addr;
  wire[2:0] prbNet_io_out_2_bits_payload_master_xact_id;
  wire[1:0] prbNet_io_out_2_bits_payload_p_type;
  wire prbNet_io_out_1_valid;
  wire[1:0] prbNet_io_out_1_bits_header_src;
  wire[1:0] prbNet_io_out_1_bits_header_dst;
  wire[25:0] prbNet_io_out_1_bits_payload_addr;
  wire[2:0] prbNet_io_out_1_bits_payload_master_xact_id;
  wire[1:0] prbNet_io_out_1_bits_payload_p_type;
  wire gntNet_io_in_0_ready;
  wire gntNet_io_out_2_valid;
  wire[1:0] gntNet_io_out_2_bits_header_src;
  wire[1:0] gntNet_io_out_2_bits_header_dst;
  wire[511:0] gntNet_io_out_2_bits_payload_data;
  wire[1:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire[2:0] gntNet_io_out_2_bits_payload_master_xact_id;
  wire[3:0] gntNet_io_out_2_bits_payload_g_type;
  wire gntNet_io_out_1_valid;
  wire[1:0] gntNet_io_out_1_bits_header_src;
  wire[1:0] gntNet_io_out_1_bits_header_dst;
  wire[511:0] gntNet_io_out_1_bits_payload_data;
  wire[1:0] gntNet_io_out_1_bits_payload_client_xact_id;
  wire[2:0] gntNet_io_out_1_bits_payload_master_xact_id;
  wire[3:0] gntNet_io_out_1_bits_payload_g_type;
  wire ackNet_io_in_2_ready;
  wire ackNet_io_in_1_ready;
  wire ackNet_io_out_0_valid;
  wire[1:0] ackNet_io_out_0_bits_header_src;
  wire[1:0] ackNet_io_out_0_bits_header_dst;
  wire[2:0] ackNet_io_out_0_bits_payload_master_xact_id;


  assign T63 = io_masters_0_finish_ready;
  assign T64 = io_clients_0_finish_bits_payload_master_xact_id;
  assign T65 = io_clients_0_finish_bits_header_dst;
  assign T66 = T67;
  assign T67 = io_clients_0_finish_bits_header_src + 2'h1;
  assign T68 = io_clients_0_finish_valid;
  assign T69 = io_clients_1_finish_bits_payload_master_xact_id;
  assign T70 = io_clients_1_finish_bits_header_dst;
  assign T71 = T72;
  assign T72 = io_clients_1_finish_bits_header_src + 2'h1;
  assign T73 = io_clients_1_finish_valid;
  assign T74 = io_clients_0_grant_ready;
  assign T75 = io_clients_1_grant_ready;
  assign T76 = io_masters_0_grant_bits_payload_g_type;
  assign T77 = io_masters_0_grant_bits_payload_master_xact_id;
  assign T78 = io_masters_0_grant_bits_payload_client_xact_id;
  assign T79 = io_masters_0_grant_bits_payload_data;
  assign T80 = T81;
  assign T81 = io_masters_0_grant_bits_header_dst + 2'h1;
  assign T82 = io_masters_0_grant_bits_header_src;
  assign T83 = io_masters_0_grant_valid;
  assign T84 = io_clients_0_probe_ready;
  assign T85 = io_clients_1_probe_ready;
  assign T86 = io_masters_0_probe_bits_payload_p_type;
  assign T87 = io_masters_0_probe_bits_payload_master_xact_id;
  assign T88 = io_masters_0_probe_bits_payload_addr;
  assign T89 = T90;
  assign T90 = io_masters_0_probe_bits_header_dst + 2'h1;
  assign T91 = io_masters_0_probe_bits_header_src;
  assign T92 = io_masters_0_probe_valid;
  assign T93 = io_masters_0_release_ready;
  assign T94 = io_clients_0_release_bits_payload_r_type;
  assign T95 = io_clients_0_release_bits_payload_data;
  assign T96 = io_clients_0_release_bits_payload_master_xact_id;
  assign T97 = io_clients_0_release_bits_payload_client_xact_id;
  assign T98 = io_clients_0_release_bits_payload_addr;
  assign T99 = io_clients_0_release_bits_header_dst;
  assign T100 = T101;
  assign T101 = io_clients_0_release_bits_header_src + 2'h1;
  assign T102 = io_clients_0_release_valid;
  assign T103 = io_clients_1_release_bits_payload_r_type;
  assign T104 = io_clients_1_release_bits_payload_data;
  assign T105 = io_clients_1_release_bits_payload_master_xact_id;
  assign T106 = io_clients_1_release_bits_payload_client_xact_id;
  assign T107 = io_clients_1_release_bits_payload_addr;
  assign T108 = io_clients_1_release_bits_header_dst;
  assign T109 = T110;
  assign T110 = io_clients_1_release_bits_header_src + 2'h1;
  assign T111 = io_clients_1_release_valid;
  assign T112 = io_masters_0_acquire_ready;
  assign T113 = io_clients_0_acquire_bits_payload_atomic_opcode;
  assign T114 = io_clients_0_acquire_bits_payload_subword_addr;
  assign T115 = io_clients_0_acquire_bits_payload_write_mask;
  assign T116 = io_clients_0_acquire_bits_payload_a_type;
  assign T117 = io_clients_0_acquire_bits_payload_data;
  assign T118 = io_clients_0_acquire_bits_payload_client_xact_id;
  assign T119 = io_clients_0_acquire_bits_payload_addr;
  assign T120 = io_clients_0_acquire_bits_header_dst;
  assign T121 = T122;
  assign T122 = io_clients_0_acquire_bits_header_src + 2'h1;
  assign T123 = io_clients_0_acquire_valid;
  assign T124 = io_clients_1_acquire_bits_payload_atomic_opcode;
  assign T125 = io_clients_1_acquire_bits_payload_subword_addr;
  assign T126 = io_clients_1_acquire_bits_payload_write_mask;
  assign T127 = io_clients_1_acquire_bits_payload_a_type;
  assign T128 = io_clients_1_acquire_bits_payload_data;
  assign T129 = io_clients_1_acquire_bits_payload_client_xact_id;
  assign T130 = io_clients_1_acquire_bits_payload_addr;
  assign T131 = io_clients_1_acquire_bits_header_dst;
  assign T132 = T133;
  assign T133 = io_clients_1_acquire_bits_header_src + 2'h1;
  assign T134 = io_clients_1_acquire_valid;
  assign io_masters_0_release_bits_payload_r_type = T0;
  assign T0 = relNet_io_out_0_bits_payload_r_type;
  assign io_masters_0_release_bits_payload_data = T1;
  assign T1 = relNet_io_out_0_bits_payload_data;
  assign io_masters_0_release_bits_payload_master_xact_id = T2;
  assign T2 = relNet_io_out_0_bits_payload_master_xact_id;
  assign io_masters_0_release_bits_payload_client_xact_id = T3;
  assign T3 = relNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_release_bits_payload_addr = T4;
  assign T4 = relNet_io_out_0_bits_payload_addr;
  assign io_masters_0_release_bits_header_dst = T5;
  assign T5 = relNet_io_out_0_bits_header_dst;
  assign io_masters_0_release_bits_header_src = T6;
  assign T6 = T7;
  assign T7 = relNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_release_valid = T8;
  assign T8 = relNet_io_out_0_valid;
  assign io_masters_0_probe_ready = T9;
  assign T9 = prbNet_io_in_0_ready;
  assign io_masters_0_finish_bits_payload_master_xact_id = T10;
  assign T10 = ackNet_io_out_0_bits_payload_master_xact_id;
  assign io_masters_0_finish_bits_header_dst = T11;
  assign T11 = ackNet_io_out_0_bits_header_dst;
  assign io_masters_0_finish_bits_header_src = T12;
  assign T12 = T13;
  assign T13 = ackNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_finish_valid = T14;
  assign T14 = ackNet_io_out_0_valid;
  assign io_masters_0_grant_ready = T15;
  assign T15 = gntNet_io_in_0_ready;
  assign io_masters_0_acquire_bits_payload_atomic_opcode = T16;
  assign T16 = acqNet_io_out_0_bits_payload_atomic_opcode;
  assign io_masters_0_acquire_bits_payload_subword_addr = T17;
  assign T17 = acqNet_io_out_0_bits_payload_subword_addr;
  assign io_masters_0_acquire_bits_payload_write_mask = T18;
  assign T18 = acqNet_io_out_0_bits_payload_write_mask;
  assign io_masters_0_acquire_bits_payload_a_type = T19;
  assign T19 = acqNet_io_out_0_bits_payload_a_type;
  assign io_masters_0_acquire_bits_payload_data = T20;
  assign T20 = acqNet_io_out_0_bits_payload_data;
  assign io_masters_0_acquire_bits_payload_client_xact_id = T21;
  assign T21 = acqNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_acquire_bits_payload_addr = T22;
  assign T22 = acqNet_io_out_0_bits_payload_addr;
  assign io_masters_0_acquire_bits_header_dst = T23;
  assign T23 = acqNet_io_out_0_bits_header_dst;
  assign io_masters_0_acquire_bits_header_src = T24;
  assign T24 = T25;
  assign T25 = acqNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_acquire_valid = T26;
  assign T26 = acqNet_io_out_0_valid;
  assign io_clients_0_release_ready = T27;
  assign T27 = relNet_io_in_1_ready;
  assign io_clients_0_probe_bits_payload_p_type = T28;
  assign T28 = prbNet_io_out_1_bits_payload_p_type;
  assign io_clients_0_probe_bits_payload_master_xact_id = T29;
  assign T29 = prbNet_io_out_1_bits_payload_master_xact_id;
  assign io_clients_0_probe_bits_payload_addr = T30;
  assign T30 = prbNet_io_out_1_bits_payload_addr;
  assign io_clients_0_probe_bits_header_dst = T31;
  assign T31 = T32;
  assign T32 = prbNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_probe_bits_header_src = T33;
  assign T33 = prbNet_io_out_1_bits_header_src;
  assign io_clients_0_probe_valid = T34;
  assign T34 = prbNet_io_out_1_valid;
  assign io_clients_0_finish_ready = T35;
  assign T35 = ackNet_io_in_1_ready;
  assign io_clients_0_grant_bits_payload_g_type = T36;
  assign T36 = gntNet_io_out_1_bits_payload_g_type;
  assign io_clients_0_grant_bits_payload_master_xact_id = T37;
  assign T37 = gntNet_io_out_1_bits_payload_master_xact_id;
  assign io_clients_0_grant_bits_payload_client_xact_id = T38;
  assign T38 = gntNet_io_out_1_bits_payload_client_xact_id;
  assign io_clients_0_grant_bits_payload_data = T39;
  assign T39 = gntNet_io_out_1_bits_payload_data;
  assign io_clients_0_grant_bits_header_dst = T40;
  assign T40 = T41;
  assign T41 = gntNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_grant_bits_header_src = T42;
  assign T42 = gntNet_io_out_1_bits_header_src;
  assign io_clients_0_grant_valid = T43;
  assign T43 = gntNet_io_out_1_valid;
  assign io_clients_0_acquire_ready = T44;
  assign T44 = acqNet_io_in_1_ready;
  assign io_clients_1_release_ready = T45;
  assign T45 = relNet_io_in_2_ready;
  assign io_clients_1_probe_bits_payload_p_type = T46;
  assign T46 = prbNet_io_out_2_bits_payload_p_type;
  assign io_clients_1_probe_bits_payload_master_xact_id = T47;
  assign T47 = prbNet_io_out_2_bits_payload_master_xact_id;
  assign io_clients_1_probe_bits_payload_addr = T48;
  assign T48 = prbNet_io_out_2_bits_payload_addr;
  assign io_clients_1_probe_bits_header_dst = T49;
  assign T49 = T50;
  assign T50 = prbNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_probe_bits_header_src = T51;
  assign T51 = prbNet_io_out_2_bits_header_src;
  assign io_clients_1_probe_valid = T52;
  assign T52 = prbNet_io_out_2_valid;
  assign io_clients_1_finish_ready = T53;
  assign T53 = ackNet_io_in_2_ready;
  assign io_clients_1_grant_bits_payload_g_type = T54;
  assign T54 = gntNet_io_out_2_bits_payload_g_type;
  assign io_clients_1_grant_bits_payload_master_xact_id = T55;
  assign T55 = gntNet_io_out_2_bits_payload_master_xact_id;
  assign io_clients_1_grant_bits_payload_client_xact_id = T56;
  assign T56 = gntNet_io_out_2_bits_payload_client_xact_id;
  assign io_clients_1_grant_bits_payload_data = T57;
  assign T57 = gntNet_io_out_2_bits_payload_data;
  assign io_clients_1_grant_bits_header_dst = T58;
  assign T58 = T59;
  assign T59 = gntNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_grant_bits_header_src = T60;
  assign T60 = gntNet_io_out_2_bits_header_src;
  assign io_clients_1_grant_valid = T61;
  assign T61 = gntNet_io_out_2_valid;
  assign io_clients_1_acquire_ready = T62;
  assign T62 = acqNet_io_in_2_ready;
  BasicCrossbar_0 acqNet(.clk(clk), .reset(reset),
       .io_in_2_ready( acqNet_io_in_2_ready ),
       .io_in_2_valid( T134 ),
       .io_in_2_bits_header_src( T132 ),
       .io_in_2_bits_header_dst( T131 ),
       .io_in_2_bits_payload_addr( T130 ),
       .io_in_2_bits_payload_client_xact_id( T129 ),
       .io_in_2_bits_payload_data( T128 ),
       .io_in_2_bits_payload_a_type( T127 ),
       .io_in_2_bits_payload_write_mask( T126 ),
       .io_in_2_bits_payload_subword_addr( T125 ),
       .io_in_2_bits_payload_atomic_opcode( T124 ),
       .io_in_1_ready( acqNet_io_in_1_ready ),
       .io_in_1_valid( T123 ),
       .io_in_1_bits_header_src( T121 ),
       .io_in_1_bits_header_dst( T120 ),
       .io_in_1_bits_payload_addr( T119 ),
       .io_in_1_bits_payload_client_xact_id( T118 ),
       .io_in_1_bits_payload_data( T117 ),
       .io_in_1_bits_payload_a_type( T116 ),
       .io_in_1_bits_payload_write_mask( T115 ),
       .io_in_1_bits_payload_subword_addr( T114 ),
       .io_in_1_bits_payload_atomic_opcode( T113 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_a_type(  )
       //.io_in_0_bits_payload_write_mask(  )
       //.io_in_0_bits_payload_subword_addr(  )
       //.io_in_0_bits_payload_atomic_opcode(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_a_type(  )
       //.io_out_2_bits_payload_write_mask(  )
       //.io_out_2_bits_payload_subword_addr(  )
       //.io_out_2_bits_payload_atomic_opcode(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_a_type(  )
       //.io_out_1_bits_payload_write_mask(  )
       //.io_out_1_bits_payload_subword_addr(  )
       //.io_out_1_bits_payload_atomic_opcode(  )
       .io_out_0_ready( T112 ),
       .io_out_0_valid( acqNet_io_out_0_valid ),
       .io_out_0_bits_header_src( acqNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( acqNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( acqNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( acqNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_data( acqNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_a_type( acqNet_io_out_0_bits_payload_a_type ),
       .io_out_0_bits_payload_write_mask( acqNet_io_out_0_bits_payload_write_mask ),
       .io_out_0_bits_payload_subword_addr( acqNet_io_out_0_bits_payload_subword_addr ),
       .io_out_0_bits_payload_atomic_opcode( acqNet_io_out_0_bits_payload_atomic_opcode )
  );
  `ifndef SYNTHESIS
    assign acqNet.io_in_0_bits_header_src = {1{$random}};
    assign acqNet.io_in_0_bits_header_dst = {1{$random}};
    assign acqNet.io_in_0_bits_payload_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign acqNet.io_in_0_bits_payload_data = {16{$random}};
    assign acqNet.io_in_0_bits_payload_a_type = {1{$random}};
    assign acqNet.io_in_0_bits_payload_write_mask = {1{$random}};
    assign acqNet.io_in_0_bits_payload_subword_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_atomic_opcode = {1{$random}};
  `endif
  BasicCrossbar_1 relNet(.clk(clk), .reset(reset),
       .io_in_2_ready( relNet_io_in_2_ready ),
       .io_in_2_valid( T111 ),
       .io_in_2_bits_header_src( T109 ),
       .io_in_2_bits_header_dst( T108 ),
       .io_in_2_bits_payload_addr( T107 ),
       .io_in_2_bits_payload_client_xact_id( T106 ),
       .io_in_2_bits_payload_master_xact_id( T105 ),
       .io_in_2_bits_payload_data( T104 ),
       .io_in_2_bits_payload_r_type( T103 ),
       .io_in_1_ready( relNet_io_in_1_ready ),
       .io_in_1_valid( T102 ),
       .io_in_1_bits_header_src( T100 ),
       .io_in_1_bits_header_dst( T99 ),
       .io_in_1_bits_payload_addr( T98 ),
       .io_in_1_bits_payload_client_xact_id( T97 ),
       .io_in_1_bits_payload_master_xact_id( T96 ),
       .io_in_1_bits_payload_data( T95 ),
       .io_in_1_bits_payload_r_type( T94 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_r_type(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_master_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_r_type(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_master_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_r_type(  )
       .io_out_0_ready( T93 ),
       .io_out_0_valid( relNet_io_out_0_valid ),
       .io_out_0_bits_header_src( relNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( relNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( relNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( relNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_master_xact_id( relNet_io_out_0_bits_payload_master_xact_id ),
       .io_out_0_bits_payload_data( relNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_r_type( relNet_io_out_0_bits_payload_r_type )
  );
  `ifndef SYNTHESIS
    assign relNet.io_in_0_bits_header_src = {1{$random}};
    assign relNet.io_in_0_bits_header_dst = {1{$random}};
    assign relNet.io_in_0_bits_payload_addr = {1{$random}};
    assign relNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_master_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_data = {16{$random}};
    assign relNet.io_in_0_bits_payload_r_type = {1{$random}};
  `endif
  BasicCrossbar_2 prbNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_addr(  )
       //.io_in_2_bits_payload_master_xact_id(  )
       //.io_in_2_bits_payload_p_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_addr(  )
       //.io_in_1_bits_payload_master_xact_id(  )
       //.io_in_1_bits_payload_p_type(  )
       .io_in_0_ready( prbNet_io_in_0_ready ),
       .io_in_0_valid( T92 ),
       .io_in_0_bits_header_src( T91 ),
       .io_in_0_bits_header_dst( T89 ),
       .io_in_0_bits_payload_addr( T88 ),
       .io_in_0_bits_payload_master_xact_id( T87 ),
       .io_in_0_bits_payload_p_type( T86 ),
       .io_out_2_ready( T85 ),
       .io_out_2_valid( prbNet_io_out_2_valid ),
       .io_out_2_bits_header_src( prbNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( prbNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_addr( prbNet_io_out_2_bits_payload_addr ),
       .io_out_2_bits_payload_master_xact_id( prbNet_io_out_2_bits_payload_master_xact_id ),
       .io_out_2_bits_payload_p_type( prbNet_io_out_2_bits_payload_p_type ),
       .io_out_1_ready( T84 ),
       .io_out_1_valid( prbNet_io_out_1_valid ),
       .io_out_1_bits_header_src( prbNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( prbNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_addr( prbNet_io_out_1_bits_payload_addr ),
       .io_out_1_bits_payload_master_xact_id( prbNet_io_out_1_bits_payload_master_xact_id ),
       .io_out_1_bits_payload_p_type( prbNet_io_out_1_bits_payload_p_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_addr(  )
       //.io_out_0_bits_payload_master_xact_id(  )
       //.io_out_0_bits_payload_p_type(  )
  );
  `ifndef SYNTHESIS
    assign prbNet.io_in_2_bits_header_src = {1{$random}};
    assign prbNet.io_in_2_bits_header_dst = {1{$random}};
    assign prbNet.io_in_2_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_2_bits_payload_master_xact_id = {1{$random}};
    assign prbNet.io_in_2_bits_payload_p_type = {1{$random}};
    assign prbNet.io_in_1_bits_header_src = {1{$random}};
    assign prbNet.io_in_1_bits_header_dst = {1{$random}};
    assign prbNet.io_in_1_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_1_bits_payload_master_xact_id = {1{$random}};
    assign prbNet.io_in_1_bits_payload_p_type = {1{$random}};
  `endif
  BasicCrossbar_3 gntNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_data(  )
       //.io_in_2_bits_payload_client_xact_id(  )
       //.io_in_2_bits_payload_master_xact_id(  )
       //.io_in_2_bits_payload_g_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_data(  )
       //.io_in_1_bits_payload_client_xact_id(  )
       //.io_in_1_bits_payload_master_xact_id(  )
       //.io_in_1_bits_payload_g_type(  )
       .io_in_0_ready( gntNet_io_in_0_ready ),
       .io_in_0_valid( T83 ),
       .io_in_0_bits_header_src( T82 ),
       .io_in_0_bits_header_dst( T80 ),
       .io_in_0_bits_payload_data( T79 ),
       .io_in_0_bits_payload_client_xact_id( T78 ),
       .io_in_0_bits_payload_master_xact_id( T77 ),
       .io_in_0_bits_payload_g_type( T76 ),
       .io_out_2_ready( T75 ),
       .io_out_2_valid( gntNet_io_out_2_valid ),
       .io_out_2_bits_header_src( gntNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( gntNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_data( gntNet_io_out_2_bits_payload_data ),
       .io_out_2_bits_payload_client_xact_id( gntNet_io_out_2_bits_payload_client_xact_id ),
       .io_out_2_bits_payload_master_xact_id( gntNet_io_out_2_bits_payload_master_xact_id ),
       .io_out_2_bits_payload_g_type( gntNet_io_out_2_bits_payload_g_type ),
       .io_out_1_ready( T74 ),
       .io_out_1_valid( gntNet_io_out_1_valid ),
       .io_out_1_bits_header_src( gntNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( gntNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_data( gntNet_io_out_1_bits_payload_data ),
       .io_out_1_bits_payload_client_xact_id( gntNet_io_out_1_bits_payload_client_xact_id ),
       .io_out_1_bits_payload_master_xact_id( gntNet_io_out_1_bits_payload_master_xact_id ),
       .io_out_1_bits_payload_g_type( gntNet_io_out_1_bits_payload_g_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_data(  )
       //.io_out_0_bits_payload_client_xact_id(  )
       //.io_out_0_bits_payload_master_xact_id(  )
       //.io_out_0_bits_payload_g_type(  )
  );
  `ifndef SYNTHESIS
    assign gntNet.io_in_2_bits_header_src = {1{$random}};
    assign gntNet.io_in_2_bits_header_dst = {1{$random}};
    assign gntNet.io_in_2_bits_payload_data = {16{$random}};
    assign gntNet.io_in_2_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_g_type = {1{$random}};
    assign gntNet.io_in_1_bits_header_src = {1{$random}};
    assign gntNet.io_in_1_bits_header_dst = {1{$random}};
    assign gntNet.io_in_1_bits_payload_data = {16{$random}};
    assign gntNet.io_in_1_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_g_type = {1{$random}};
  `endif
  BasicCrossbar_4 ackNet(.clk(clk), .reset(reset),
       .io_in_2_ready( ackNet_io_in_2_ready ),
       .io_in_2_valid( T73 ),
       .io_in_2_bits_header_src( T71 ),
       .io_in_2_bits_header_dst( T70 ),
       .io_in_2_bits_payload_master_xact_id( T69 ),
       .io_in_1_ready( ackNet_io_in_1_ready ),
       .io_in_1_valid( T68 ),
       .io_in_1_bits_header_src( T66 ),
       .io_in_1_bits_header_dst( T65 ),
       .io_in_1_bits_payload_master_xact_id( T64 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_master_xact_id(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_master_xact_id(  )
       .io_out_0_ready( T63 ),
       .io_out_0_valid( ackNet_io_out_0_valid ),
       .io_out_0_bits_header_src( ackNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( ackNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_master_xact_id( ackNet_io_out_0_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign ackNet.io_in_0_bits_header_src = {1{$random}};
    assign ackNet.io_in_0_bits_header_dst = {1{$random}};
    assign ackNet.io_in_0_bits_payload_master_xact_id = {1{$random}};
  `endif
endmodule

module VoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[1:0] io_inner_probe_bits_header_src
    //output[1:0] io_inner_probe_bits_header_dst
    //output[25:0] io_inner_probe_bits_payload_addr
    //output[2:0] io_inner_probe_bits_payload_master_xact_id
    //output[1:0] io_inner_probe_bits_payload_p_type
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [1:0] state;
  wire[1:0] T38;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg [25:0] xact_addr;
  wire[25:0] T20;
  wire[3:0] T21;
  wire[2:0] T22;
  wire[5:0] T23;
  wire[2:0] T24;
  wire[511:0] T25;
  reg [511:0] xact_data;
  wire[511:0] T26;
  wire[1:0] T27;
  wire[25:0] T28;
  wire[3:0] T29;
  wire[3:0] T30;
  wire T31;
  reg [2:0] xact_r_type;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[1:0] T34;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T35;
  wire[511:0] T36;
  wire[1:0] T39;
  reg  init_client_id;
  wire T40;
  wire[1:0] T41;
  wire[1:0] T37;
  wire[1:0] T42;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    xact_r_type = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T19 & T1;
  assign T1 = state != 2'h0;
  assign T38 = reset ? 2'h0 : T2;
  assign T2 = T17 ? 2'h0 : T3;
  assign T3 = T15 ? 2'h2 : T4;
  assign T4 = T13 ? T5 : state;
  assign T5 = T6 ? 2'h1 : 2'h2;
  assign T6 = T8 | T7;
  assign T7 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T8 = T10 | T9;
  assign T9 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T10 = T12 | T11;
  assign T11 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T12 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T13 = T14 & io_inner_release_valid;
  assign T14 = 2'h0 == state;
  assign T15 = T16 & io_outer_acquire_ready;
  assign T16 = 2'h1 == state;
  assign T17 = T18 & io_inner_grant_ready;
  assign T18 = 2'h2 == state;
  assign T19 = xact_addr == io_inner_release_bits_payload_addr;
  assign T20 = T13 ? io_inner_release_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = 1'h0;
  assign io_outer_grant_ready = 1'h0;
  assign io_outer_acquire_bits_payload_atomic_opcode = T21;
  assign T21 = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T22;
  assign T22 = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T23;
  assign T23 = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T24;
  assign T24 = 3'h3;
  assign io_outer_acquire_bits_payload_data = T25;
  assign T25 = xact_data;
  assign T26 = T13 ? io_inner_release_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T27;
  assign T27 = 2'h0;
  assign io_outer_acquire_bits_payload_addr = T28;
  assign T28 = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T16;
  assign io_inner_release_ready = T14;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_grant_bits_payload_g_type = T29;
  assign T29 = T30;
  assign T30 = T31 ? 4'h0 : 4'h3;
  assign T31 = xact_r_type == 3'h0;
  assign T32 = T13 ? io_inner_release_bits_payload_r_type : xact_r_type;
  assign io_inner_grant_bits_payload_master_xact_id = T33;
  assign T33 = 3'h0;
  assign io_inner_grant_bits_payload_client_xact_id = T34;
  assign T34 = xact_client_xact_id;
  assign T35 = T13 ? io_inner_release_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T36;
  assign T36 = 512'h0;
  assign io_inner_grant_bits_header_dst = T39;
  assign T39 = {1'h0, init_client_id};
  assign T40 = T41[1'h0:1'h0];
  assign T41 = reset ? 2'h0 : T37;
  assign T37 = T13 ? io_inner_release_bits_header_src : T42;
  assign T42 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T18;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T17) begin
      state <= 2'h0;
    end else if(T15) begin
      state <= 2'h2;
    end else if(T13) begin
      state <= T5;
    end
    if(T13) begin
      xact_addr <= io_inner_release_bits_payload_addr;
    end
    if(T13) begin
      xact_data <= io_inner_release_bits_payload_data;
    end
    if(T13) begin
      xact_r_type <= io_inner_release_bits_payload_r_type;
    end
    if(T13) begin
      xact_client_xact_id <= io_inner_release_bits_payload_client_xact_id;
    end
    init_client_id <= T40;
  end
endmodule

module AcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T154;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T155;
  wire[1:0] T156;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T157;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T158;
  wire T38;
  wire[1:0] T159;
  wire T39;
  wire[1:0] T160;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[3:0] T72;
  wire T73;
  reg  init_sharer_cnt;
  wire T161;
  wire[1:0] T162;
  wire[1:0] T74;
  wire[1:0] T163;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire[2:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg [25:0] xact_addr;
  wire[25:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T97;
  wire[2:0] T98;
  wire[2:0] T99;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T100;
  wire[5:0] T101;
  wire[5:0] T102;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T103;
  wire[2:0] T104;
  wire[2:0] T105;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T106;
  wire[511:0] T107;
  wire[511:0] T108;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T113;
  wire[25:0] T114;
  wire[25:0] T115;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T116;
  wire T117;
  wire T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[25:0] T135;
  wire[1:0] T164;
  wire T165;
  wire T166;
  reg [1:0] probe_flags;
  wire[1:0] T167;
  wire[1:0] T136;
  wire[1:0] T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire[3:0] T144;
  wire[2:0] T145;
  wire[1:0] T146;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T147;
  wire[511:0] T148;
  wire[1:0] T168;
  reg  init_client_id;
  wire T169;
  wire[1:0] T170;
  wire[1:0] T149;
  wire[1:0] T171;
  wire T150;
  wire T151;
  wire T152;
  wire T153;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T154 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T81 : T4;
  assign T4 = T79 ? T78 : T5;
  assign T5 = T76 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T155 = T156[1'h0:1'h0];
  assign T156 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T160 : T33;
  assign T33 = T52 ? T159 : T34;
  assign T34 = T21 ? T35 : T157;
  assign T157 = {1'h0, release_count};
  assign T35 = T158 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T158 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T159 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T160 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T75 ? T72 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = T73 ? 4'h1 : 4'h2;
  assign T73 = 1'h0 < init_sharer_cnt;
  assign T161 = T162[1'h0:1'h0];
  assign T162 = reset ? 2'h0 : T74;
  assign T74 = T21 ? 2'h2 : T163;
  assign T163 = {1'h0, init_sharer_cnt};
  assign T75 = xact_a_type == 3'h0;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h2 == state;
  assign T78 = pending_outer_read ? 3'h2 : 3'h4;
  assign T79 = T80 & io_outer_acquire_ready;
  assign T80 = 3'h3 == state;
  assign T81 = T82 ? 3'h5 : 3'h0;
  assign T82 = grant_type != 4'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_master_xact_id == 3'h1;
  assign T88 = 3'h5 == state;
  assign T89 = xact_addr == io_inner_release_bits_payload_addr;
  assign T90 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T91;
  assign T91 = T93 & T92;
  assign T92 = state != 3'h0;
  assign T93 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T94;
  assign T94 = T80 ? outer_write_acq_atomic_opcode : T95;
  assign T95 = T77 ? outer_read_atomic_opcode : T96;
  assign T96 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T97;
  assign T97 = T80 ? outer_write_acq_subword_addr : T98;
  assign T98 = T77 ? outer_read_subword_addr : T99;
  assign T99 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T100;
  assign T100 = T80 ? outer_write_acq_write_mask : T101;
  assign T101 = T77 ? outer_read_write_mask : T102;
  assign T102 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T103;
  assign T103 = T80 ? outer_write_acq_a_type : T104;
  assign T104 = T77 ? outer_read_a_type : T105;
  assign T105 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T106;
  assign T106 = T80 ? outer_write_acq_data : T107;
  assign T107 = T77 ? outer_read_data : T108;
  assign T108 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T109 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T110;
  assign T110 = T80 ? outer_write_acq_client_xact_id : T111;
  assign T111 = T77 ? outer_read_client_xact_id : T112;
  assign T112 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 2'h1;
  assign outer_read_client_xact_id = 2'h1;
  assign outer_write_acq_client_xact_id = 2'h1;
  assign io_outer_acquire_bits_payload_addr = T113;
  assign T113 = T80 ? outer_write_acq_addr : T114;
  assign T114 = T77 ? outer_read_addr : T115;
  assign T115 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T116;
  assign T116 = T80 ? 1'h1 : T117;
  assign T117 = T77 ? 1'h1 : T53;
  assign io_inner_release_ready = T118;
  assign T118 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T119;
  assign T119 = T120;
  assign T120 = T133 ? 2'h1 : T121;
  assign T121 = T132 ? 2'h0 : T122;
  assign T122 = T131 ? 2'h2 : T123;
  assign T123 = T130 ? 2'h0 : T124;
  assign T124 = T129 ? 2'h2 : T125;
  assign T125 = T128 ? 2'h0 : T126;
  assign T126 = T127 ? 2'h0 : 2'h2;
  assign T127 = xact_a_type == 3'h6;
  assign T128 = xact_a_type == 3'h5;
  assign T129 = xact_a_type == 3'h4;
  assign T130 = xact_a_type == 3'h3;
  assign T131 = xact_a_type == 3'h2;
  assign T132 = xact_a_type == 3'h1;
  assign T133 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T134;
  assign T134 = 3'h1;
  assign io_inner_probe_bits_payload_addr = T135;
  assign T135 = xact_addr;
  assign io_inner_probe_bits_header_dst = T164;
  assign T164 = {1'h0, T165};
  assign T165 = T166 == 1'h0;
  assign T166 = probe_flags[1'h0:1'h0];
  assign T167 = reset ? 2'h0 : T136;
  assign T136 = T141 ? T138 : T137;
  assign T137 = T21 ? probe_initial_flags : probe_flags;
  assign T138 = probe_flags & T139;
  assign T139 = ~ T140;
  assign T140 = 1'h1 << T165;
  assign T141 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T142;
  assign T142 = T51 ? T143 : 1'h0;
  assign T143 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T144;
  assign T144 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T145;
  assign T145 = 3'h1;
  assign io_inner_grant_bits_payload_client_xact_id = T146;
  assign T146 = xact_client_xact_id;
  assign T147 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T148;
  assign T148 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T168;
  assign T168 = {1'h0, init_client_id};
  assign T169 = T170[1'h0:1'h0];
  assign T170 = reset ? 2'h0 : T149;
  assign T149 = T21 ? io_inner_acquire_bits_header_src : T171;
  assign T171 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T150;
  assign T150 = T151 ? 1'h1 : T84;
  assign T151 = T88 & T152;
  assign T152 = io_outer_grant_valid & T153;
  assign T153 = io_outer_grant_bits_payload_client_xact_id == 2'h1;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T81;
    end else if(T79) begin
      state <= T78;
    end else if(T76) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T155;
    init_sharer_cnt <= T161;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T141) begin
      probe_flags <= T138;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T169;
  end
endmodule

module AcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T154;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T155;
  wire[1:0] T156;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T157;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T158;
  wire T38;
  wire[1:0] T159;
  wire T39;
  wire[1:0] T160;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[3:0] T72;
  wire T73;
  reg  init_sharer_cnt;
  wire T161;
  wire[1:0] T162;
  wire[1:0] T74;
  wire[1:0] T163;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire[2:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg [25:0] xact_addr;
  wire[25:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T97;
  wire[2:0] T98;
  wire[2:0] T99;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T100;
  wire[5:0] T101;
  wire[5:0] T102;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T103;
  wire[2:0] T104;
  wire[2:0] T105;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T106;
  wire[511:0] T107;
  wire[511:0] T108;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T113;
  wire[25:0] T114;
  wire[25:0] T115;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T116;
  wire T117;
  wire T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[25:0] T135;
  wire[1:0] T164;
  wire T165;
  wire T166;
  reg [1:0] probe_flags;
  wire[1:0] T167;
  wire[1:0] T136;
  wire[1:0] T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire[3:0] T144;
  wire[2:0] T145;
  wire[1:0] T146;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T147;
  wire[511:0] T148;
  wire[1:0] T168;
  reg  init_client_id;
  wire T169;
  wire[1:0] T170;
  wire[1:0] T149;
  wire[1:0] T171;
  wire T150;
  wire T151;
  wire T152;
  wire T153;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T154 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T81 : T4;
  assign T4 = T79 ? T78 : T5;
  assign T5 = T76 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T155 = T156[1'h0:1'h0];
  assign T156 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T160 : T33;
  assign T33 = T52 ? T159 : T34;
  assign T34 = T21 ? T35 : T157;
  assign T157 = {1'h0, release_count};
  assign T35 = T158 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T158 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T159 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T160 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T75 ? T72 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = T73 ? 4'h1 : 4'h2;
  assign T73 = 1'h0 < init_sharer_cnt;
  assign T161 = T162[1'h0:1'h0];
  assign T162 = reset ? 2'h0 : T74;
  assign T74 = T21 ? 2'h2 : T163;
  assign T163 = {1'h0, init_sharer_cnt};
  assign T75 = xact_a_type == 3'h0;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h2 == state;
  assign T78 = pending_outer_read ? 3'h2 : 3'h4;
  assign T79 = T80 & io_outer_acquire_ready;
  assign T80 = 3'h3 == state;
  assign T81 = T82 ? 3'h5 : 3'h0;
  assign T82 = grant_type != 4'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_master_xact_id == 3'h2;
  assign T88 = 3'h5 == state;
  assign T89 = xact_addr == io_inner_release_bits_payload_addr;
  assign T90 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T91;
  assign T91 = T93 & T92;
  assign T92 = state != 3'h0;
  assign T93 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T94;
  assign T94 = T80 ? outer_write_acq_atomic_opcode : T95;
  assign T95 = T77 ? outer_read_atomic_opcode : T96;
  assign T96 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T97;
  assign T97 = T80 ? outer_write_acq_subword_addr : T98;
  assign T98 = T77 ? outer_read_subword_addr : T99;
  assign T99 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T100;
  assign T100 = T80 ? outer_write_acq_write_mask : T101;
  assign T101 = T77 ? outer_read_write_mask : T102;
  assign T102 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T103;
  assign T103 = T80 ? outer_write_acq_a_type : T104;
  assign T104 = T77 ? outer_read_a_type : T105;
  assign T105 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T106;
  assign T106 = T80 ? outer_write_acq_data : T107;
  assign T107 = T77 ? outer_read_data : T108;
  assign T108 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T109 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T110;
  assign T110 = T80 ? outer_write_acq_client_xact_id : T111;
  assign T111 = T77 ? outer_read_client_xact_id : T112;
  assign T112 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 2'h2;
  assign outer_read_client_xact_id = 2'h2;
  assign outer_write_acq_client_xact_id = 2'h2;
  assign io_outer_acquire_bits_payload_addr = T113;
  assign T113 = T80 ? outer_write_acq_addr : T114;
  assign T114 = T77 ? outer_read_addr : T115;
  assign T115 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T116;
  assign T116 = T80 ? 1'h1 : T117;
  assign T117 = T77 ? 1'h1 : T53;
  assign io_inner_release_ready = T118;
  assign T118 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T119;
  assign T119 = T120;
  assign T120 = T133 ? 2'h1 : T121;
  assign T121 = T132 ? 2'h0 : T122;
  assign T122 = T131 ? 2'h2 : T123;
  assign T123 = T130 ? 2'h0 : T124;
  assign T124 = T129 ? 2'h2 : T125;
  assign T125 = T128 ? 2'h0 : T126;
  assign T126 = T127 ? 2'h0 : 2'h2;
  assign T127 = xact_a_type == 3'h6;
  assign T128 = xact_a_type == 3'h5;
  assign T129 = xact_a_type == 3'h4;
  assign T130 = xact_a_type == 3'h3;
  assign T131 = xact_a_type == 3'h2;
  assign T132 = xact_a_type == 3'h1;
  assign T133 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T134;
  assign T134 = 3'h2;
  assign io_inner_probe_bits_payload_addr = T135;
  assign T135 = xact_addr;
  assign io_inner_probe_bits_header_dst = T164;
  assign T164 = {1'h0, T165};
  assign T165 = T166 == 1'h0;
  assign T166 = probe_flags[1'h0:1'h0];
  assign T167 = reset ? 2'h0 : T136;
  assign T136 = T141 ? T138 : T137;
  assign T137 = T21 ? probe_initial_flags : probe_flags;
  assign T138 = probe_flags & T139;
  assign T139 = ~ T140;
  assign T140 = 1'h1 << T165;
  assign T141 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T142;
  assign T142 = T51 ? T143 : 1'h0;
  assign T143 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T144;
  assign T144 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T145;
  assign T145 = 3'h2;
  assign io_inner_grant_bits_payload_client_xact_id = T146;
  assign T146 = xact_client_xact_id;
  assign T147 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T148;
  assign T148 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T168;
  assign T168 = {1'h0, init_client_id};
  assign T169 = T170[1'h0:1'h0];
  assign T170 = reset ? 2'h0 : T149;
  assign T149 = T21 ? io_inner_acquire_bits_header_src : T171;
  assign T171 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T150;
  assign T150 = T151 ? 1'h1 : T84;
  assign T151 = T88 & T152;
  assign T152 = io_outer_grant_valid & T153;
  assign T153 = io_outer_grant_bits_payload_client_xact_id == 2'h2;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T81;
    end else if(T79) begin
      state <= T78;
    end else if(T76) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T155;
    init_sharer_cnt <= T161;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T141) begin
      probe_flags <= T138;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T169;
  end
endmodule

module AcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T154;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T155;
  wire[1:0] T156;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T157;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T158;
  wire T38;
  wire[1:0] T159;
  wire T39;
  wire[1:0] T160;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[3:0] T72;
  wire T73;
  reg  init_sharer_cnt;
  wire T161;
  wire[1:0] T162;
  wire[1:0] T74;
  wire[1:0] T163;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire[2:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg [25:0] xact_addr;
  wire[25:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T97;
  wire[2:0] T98;
  wire[2:0] T99;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T100;
  wire[5:0] T101;
  wire[5:0] T102;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T103;
  wire[2:0] T104;
  wire[2:0] T105;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T106;
  wire[511:0] T107;
  wire[511:0] T108;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T113;
  wire[25:0] T114;
  wire[25:0] T115;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T116;
  wire T117;
  wire T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[25:0] T135;
  wire[1:0] T164;
  wire T165;
  wire T166;
  reg [1:0] probe_flags;
  wire[1:0] T167;
  wire[1:0] T136;
  wire[1:0] T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire[3:0] T144;
  wire[2:0] T145;
  wire[1:0] T146;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T147;
  wire[511:0] T148;
  wire[1:0] T168;
  reg  init_client_id;
  wire T169;
  wire[1:0] T170;
  wire[1:0] T149;
  wire[1:0] T171;
  wire T150;
  wire T151;
  wire T152;
  wire T153;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T154 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T81 : T4;
  assign T4 = T79 ? T78 : T5;
  assign T5 = T76 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T155 = T156[1'h0:1'h0];
  assign T156 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T160 : T33;
  assign T33 = T52 ? T159 : T34;
  assign T34 = T21 ? T35 : T157;
  assign T157 = {1'h0, release_count};
  assign T35 = T158 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T158 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T159 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T160 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T75 ? T72 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = T73 ? 4'h1 : 4'h2;
  assign T73 = 1'h0 < init_sharer_cnt;
  assign T161 = T162[1'h0:1'h0];
  assign T162 = reset ? 2'h0 : T74;
  assign T74 = T21 ? 2'h2 : T163;
  assign T163 = {1'h0, init_sharer_cnt};
  assign T75 = xact_a_type == 3'h0;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h2 == state;
  assign T78 = pending_outer_read ? 3'h2 : 3'h4;
  assign T79 = T80 & io_outer_acquire_ready;
  assign T80 = 3'h3 == state;
  assign T81 = T82 ? 3'h5 : 3'h0;
  assign T82 = grant_type != 4'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_master_xact_id == 3'h3;
  assign T88 = 3'h5 == state;
  assign T89 = xact_addr == io_inner_release_bits_payload_addr;
  assign T90 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T91;
  assign T91 = T93 & T92;
  assign T92 = state != 3'h0;
  assign T93 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T94;
  assign T94 = T80 ? outer_write_acq_atomic_opcode : T95;
  assign T95 = T77 ? outer_read_atomic_opcode : T96;
  assign T96 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T97;
  assign T97 = T80 ? outer_write_acq_subword_addr : T98;
  assign T98 = T77 ? outer_read_subword_addr : T99;
  assign T99 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T100;
  assign T100 = T80 ? outer_write_acq_write_mask : T101;
  assign T101 = T77 ? outer_read_write_mask : T102;
  assign T102 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T103;
  assign T103 = T80 ? outer_write_acq_a_type : T104;
  assign T104 = T77 ? outer_read_a_type : T105;
  assign T105 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T106;
  assign T106 = T80 ? outer_write_acq_data : T107;
  assign T107 = T77 ? outer_read_data : T108;
  assign T108 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T109 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T110;
  assign T110 = T80 ? outer_write_acq_client_xact_id : T111;
  assign T111 = T77 ? outer_read_client_xact_id : T112;
  assign T112 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 2'h3;
  assign outer_read_client_xact_id = 2'h3;
  assign outer_write_acq_client_xact_id = 2'h3;
  assign io_outer_acquire_bits_payload_addr = T113;
  assign T113 = T80 ? outer_write_acq_addr : T114;
  assign T114 = T77 ? outer_read_addr : T115;
  assign T115 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T116;
  assign T116 = T80 ? 1'h1 : T117;
  assign T117 = T77 ? 1'h1 : T53;
  assign io_inner_release_ready = T118;
  assign T118 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T119;
  assign T119 = T120;
  assign T120 = T133 ? 2'h1 : T121;
  assign T121 = T132 ? 2'h0 : T122;
  assign T122 = T131 ? 2'h2 : T123;
  assign T123 = T130 ? 2'h0 : T124;
  assign T124 = T129 ? 2'h2 : T125;
  assign T125 = T128 ? 2'h0 : T126;
  assign T126 = T127 ? 2'h0 : 2'h2;
  assign T127 = xact_a_type == 3'h6;
  assign T128 = xact_a_type == 3'h5;
  assign T129 = xact_a_type == 3'h4;
  assign T130 = xact_a_type == 3'h3;
  assign T131 = xact_a_type == 3'h2;
  assign T132 = xact_a_type == 3'h1;
  assign T133 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T134;
  assign T134 = 3'h3;
  assign io_inner_probe_bits_payload_addr = T135;
  assign T135 = xact_addr;
  assign io_inner_probe_bits_header_dst = T164;
  assign T164 = {1'h0, T165};
  assign T165 = T166 == 1'h0;
  assign T166 = probe_flags[1'h0:1'h0];
  assign T167 = reset ? 2'h0 : T136;
  assign T136 = T141 ? T138 : T137;
  assign T137 = T21 ? probe_initial_flags : probe_flags;
  assign T138 = probe_flags & T139;
  assign T139 = ~ T140;
  assign T140 = 1'h1 << T165;
  assign T141 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T142;
  assign T142 = T51 ? T143 : 1'h0;
  assign T143 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T144;
  assign T144 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T145;
  assign T145 = 3'h3;
  assign io_inner_grant_bits_payload_client_xact_id = T146;
  assign T146 = xact_client_xact_id;
  assign T147 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T148;
  assign T148 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T168;
  assign T168 = {1'h0, init_client_id};
  assign T169 = T170[1'h0:1'h0];
  assign T170 = reset ? 2'h0 : T149;
  assign T149 = T21 ? io_inner_acquire_bits_header_src : T171;
  assign T171 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T150;
  assign T150 = T151 ? 1'h1 : T84;
  assign T151 = T88 & T152;
  assign T152 = io_outer_grant_valid & T153;
  assign T153 = io_outer_grant_bits_payload_client_xact_id == 2'h3;
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T81;
    end else if(T79) begin
      state <= T78;
    end else if(T76) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T155;
    init_sharer_cnt <= T161;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T141) begin
      probe_flags <= T138;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T169;
  end
endmodule

module AcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T154;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T155;
  wire[1:0] T156;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T157;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T158;
  wire T38;
  wire[1:0] T159;
  wire T39;
  wire[1:0] T160;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[3:0] T72;
  wire T73;
  reg  init_sharer_cnt;
  wire T161;
  wire[1:0] T162;
  wire[1:0] T74;
  wire[1:0] T163;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire[2:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg [25:0] xact_addr;
  wire[25:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T97;
  wire[2:0] T98;
  wire[2:0] T99;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T100;
  wire[5:0] T101;
  wire[5:0] T102;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T103;
  wire[2:0] T104;
  wire[2:0] T105;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T106;
  wire[511:0] T107;
  wire[511:0] T108;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T113;
  wire[25:0] T114;
  wire[25:0] T115;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T116;
  wire T117;
  wire T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[25:0] T135;
  wire[1:0] T164;
  wire T165;
  wire T166;
  reg [1:0] probe_flags;
  wire[1:0] T167;
  wire[1:0] T136;
  wire[1:0] T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire[3:0] T144;
  wire[2:0] T145;
  wire[1:0] T146;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T147;
  wire[511:0] T148;
  wire[1:0] T168;
  reg  init_client_id;
  wire T169;
  wire[1:0] T170;
  wire[1:0] T149;
  wire[1:0] T171;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire[2:0] T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T154 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T81 : T4;
  assign T4 = T79 ? T78 : T5;
  assign T5 = T76 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T155 = T156[1'h0:1'h0];
  assign T156 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T160 : T33;
  assign T33 = T52 ? T159 : T34;
  assign T34 = T21 ? T35 : T157;
  assign T157 = {1'h0, release_count};
  assign T35 = T158 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T158 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T159 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T160 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T75 ? T72 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = T73 ? 4'h1 : 4'h2;
  assign T73 = 1'h0 < init_sharer_cnt;
  assign T161 = T162[1'h0:1'h0];
  assign T162 = reset ? 2'h0 : T74;
  assign T74 = T21 ? 2'h2 : T163;
  assign T163 = {1'h0, init_sharer_cnt};
  assign T75 = xact_a_type == 3'h0;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h2 == state;
  assign T78 = pending_outer_read ? 3'h2 : 3'h4;
  assign T79 = T80 & io_outer_acquire_ready;
  assign T80 = 3'h3 == state;
  assign T81 = T82 ? 3'h5 : 3'h0;
  assign T82 = grant_type != 4'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_master_xact_id == 3'h4;
  assign T88 = 3'h5 == state;
  assign T89 = xact_addr == io_inner_release_bits_payload_addr;
  assign T90 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T91;
  assign T91 = T93 & T92;
  assign T92 = state != 3'h0;
  assign T93 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T94;
  assign T94 = T80 ? outer_write_acq_atomic_opcode : T95;
  assign T95 = T77 ? outer_read_atomic_opcode : T96;
  assign T96 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T97;
  assign T97 = T80 ? outer_write_acq_subword_addr : T98;
  assign T98 = T77 ? outer_read_subword_addr : T99;
  assign T99 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T100;
  assign T100 = T80 ? outer_write_acq_write_mask : T101;
  assign T101 = T77 ? outer_read_write_mask : T102;
  assign T102 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T103;
  assign T103 = T80 ? outer_write_acq_a_type : T104;
  assign T104 = T77 ? outer_read_a_type : T105;
  assign T105 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T106;
  assign T106 = T80 ? outer_write_acq_data : T107;
  assign T107 = T77 ? outer_read_data : T108;
  assign T108 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T109 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T110;
  assign T110 = T80 ? outer_write_acq_client_xact_id : T111;
  assign T111 = T77 ? outer_read_client_xact_id : T112;
  assign T112 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 2'h0;
  assign outer_read_client_xact_id = 2'h0;
  assign outer_write_acq_client_xact_id = 2'h0;
  assign io_outer_acquire_bits_payload_addr = T113;
  assign T113 = T80 ? outer_write_acq_addr : T114;
  assign T114 = T77 ? outer_read_addr : T115;
  assign T115 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T116;
  assign T116 = T80 ? 1'h1 : T117;
  assign T117 = T77 ? 1'h1 : T53;
  assign io_inner_release_ready = T118;
  assign T118 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T119;
  assign T119 = T120;
  assign T120 = T133 ? 2'h1 : T121;
  assign T121 = T132 ? 2'h0 : T122;
  assign T122 = T131 ? 2'h2 : T123;
  assign T123 = T130 ? 2'h0 : T124;
  assign T124 = T129 ? 2'h2 : T125;
  assign T125 = T128 ? 2'h0 : T126;
  assign T126 = T127 ? 2'h0 : 2'h2;
  assign T127 = xact_a_type == 3'h6;
  assign T128 = xact_a_type == 3'h5;
  assign T129 = xact_a_type == 3'h4;
  assign T130 = xact_a_type == 3'h3;
  assign T131 = xact_a_type == 3'h2;
  assign T132 = xact_a_type == 3'h1;
  assign T133 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T134;
  assign T134 = 3'h4;
  assign io_inner_probe_bits_payload_addr = T135;
  assign T135 = xact_addr;
  assign io_inner_probe_bits_header_dst = T164;
  assign T164 = {1'h0, T165};
  assign T165 = T166 == 1'h0;
  assign T166 = probe_flags[1'h0:1'h0];
  assign T167 = reset ? 2'h0 : T136;
  assign T136 = T141 ? T138 : T137;
  assign T137 = T21 ? probe_initial_flags : probe_flags;
  assign T138 = probe_flags & T139;
  assign T139 = ~ T140;
  assign T140 = 1'h1 << T165;
  assign T141 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T142;
  assign T142 = T51 ? T143 : 1'h0;
  assign T143 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T144;
  assign T144 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T145;
  assign T145 = 3'h4;
  assign io_inner_grant_bits_payload_client_xact_id = T146;
  assign T146 = xact_client_xact_id;
  assign T147 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T148;
  assign T148 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T168;
  assign T168 = {1'h0, init_client_id};
  assign T169 = T170[1'h0:1'h0];
  assign T170 = reset ? 2'h0 : T149;
  assign T149 = T21 ? io_inner_acquire_bits_header_src : T171;
  assign T171 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T150;
  assign T150 = T151 ? 1'h1 : T84;
  assign T151 = T88 & T152;
  assign T152 = io_outer_grant_valid & T153;
  assign T153 = T172 == 3'h4;
  assign T172 = {1'h0, io_outer_grant_bits_payload_client_xact_id};
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T81;
    end else if(T79) begin
      state <= T78;
    end else if(T76) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T155;
    init_sharer_cnt <= T161;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T141) begin
      probe_flags <= T138;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T169;
  end
endmodule

module AcquireTracker_4(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T154;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T155;
  wire[1:0] T156;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T157;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T158;
  wire T38;
  wire[1:0] T159;
  wire T39;
  wire[1:0] T160;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[3:0] T72;
  wire T73;
  reg  init_sharer_cnt;
  wire T161;
  wire[1:0] T162;
  wire[1:0] T74;
  wire[1:0] T163;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire[2:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg [25:0] xact_addr;
  wire[25:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T97;
  wire[2:0] T98;
  wire[2:0] T99;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T100;
  wire[5:0] T101;
  wire[5:0] T102;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T103;
  wire[2:0] T104;
  wire[2:0] T105;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T106;
  wire[511:0] T107;
  wire[511:0] T108;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T113;
  wire[25:0] T114;
  wire[25:0] T115;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T116;
  wire T117;
  wire T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[25:0] T135;
  wire[1:0] T164;
  wire T165;
  wire T166;
  reg [1:0] probe_flags;
  wire[1:0] T167;
  wire[1:0] T136;
  wire[1:0] T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire[3:0] T144;
  wire[2:0] T145;
  wire[1:0] T146;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T147;
  wire[511:0] T148;
  wire[1:0] T168;
  reg  init_client_id;
  wire T169;
  wire[1:0] T170;
  wire[1:0] T149;
  wire[1:0] T171;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire[2:0] T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T154 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T81 : T4;
  assign T4 = T79 ? T78 : T5;
  assign T5 = T76 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T155 = T156[1'h0:1'h0];
  assign T156 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T160 : T33;
  assign T33 = T52 ? T159 : T34;
  assign T34 = T21 ? T35 : T157;
  assign T157 = {1'h0, release_count};
  assign T35 = T158 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T158 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T159 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T160 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T75 ? T72 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = T73 ? 4'h1 : 4'h2;
  assign T73 = 1'h0 < init_sharer_cnt;
  assign T161 = T162[1'h0:1'h0];
  assign T162 = reset ? 2'h0 : T74;
  assign T74 = T21 ? 2'h2 : T163;
  assign T163 = {1'h0, init_sharer_cnt};
  assign T75 = xact_a_type == 3'h0;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h2 == state;
  assign T78 = pending_outer_read ? 3'h2 : 3'h4;
  assign T79 = T80 & io_outer_acquire_ready;
  assign T80 = 3'h3 == state;
  assign T81 = T82 ? 3'h5 : 3'h0;
  assign T82 = grant_type != 4'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_master_xact_id == 3'h5;
  assign T88 = 3'h5 == state;
  assign T89 = xact_addr == io_inner_release_bits_payload_addr;
  assign T90 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T91;
  assign T91 = T93 & T92;
  assign T92 = state != 3'h0;
  assign T93 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T94;
  assign T94 = T80 ? outer_write_acq_atomic_opcode : T95;
  assign T95 = T77 ? outer_read_atomic_opcode : T96;
  assign T96 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T97;
  assign T97 = T80 ? outer_write_acq_subword_addr : T98;
  assign T98 = T77 ? outer_read_subword_addr : T99;
  assign T99 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T100;
  assign T100 = T80 ? outer_write_acq_write_mask : T101;
  assign T101 = T77 ? outer_read_write_mask : T102;
  assign T102 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T103;
  assign T103 = T80 ? outer_write_acq_a_type : T104;
  assign T104 = T77 ? outer_read_a_type : T105;
  assign T105 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T106;
  assign T106 = T80 ? outer_write_acq_data : T107;
  assign T107 = T77 ? outer_read_data : T108;
  assign T108 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T109 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T110;
  assign T110 = T80 ? outer_write_acq_client_xact_id : T111;
  assign T111 = T77 ? outer_read_client_xact_id : T112;
  assign T112 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 2'h1;
  assign outer_read_client_xact_id = 2'h1;
  assign outer_write_acq_client_xact_id = 2'h1;
  assign io_outer_acquire_bits_payload_addr = T113;
  assign T113 = T80 ? outer_write_acq_addr : T114;
  assign T114 = T77 ? outer_read_addr : T115;
  assign T115 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T116;
  assign T116 = T80 ? 1'h1 : T117;
  assign T117 = T77 ? 1'h1 : T53;
  assign io_inner_release_ready = T118;
  assign T118 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T119;
  assign T119 = T120;
  assign T120 = T133 ? 2'h1 : T121;
  assign T121 = T132 ? 2'h0 : T122;
  assign T122 = T131 ? 2'h2 : T123;
  assign T123 = T130 ? 2'h0 : T124;
  assign T124 = T129 ? 2'h2 : T125;
  assign T125 = T128 ? 2'h0 : T126;
  assign T126 = T127 ? 2'h0 : 2'h2;
  assign T127 = xact_a_type == 3'h6;
  assign T128 = xact_a_type == 3'h5;
  assign T129 = xact_a_type == 3'h4;
  assign T130 = xact_a_type == 3'h3;
  assign T131 = xact_a_type == 3'h2;
  assign T132 = xact_a_type == 3'h1;
  assign T133 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T134;
  assign T134 = 3'h5;
  assign io_inner_probe_bits_payload_addr = T135;
  assign T135 = xact_addr;
  assign io_inner_probe_bits_header_dst = T164;
  assign T164 = {1'h0, T165};
  assign T165 = T166 == 1'h0;
  assign T166 = probe_flags[1'h0:1'h0];
  assign T167 = reset ? 2'h0 : T136;
  assign T136 = T141 ? T138 : T137;
  assign T137 = T21 ? probe_initial_flags : probe_flags;
  assign T138 = probe_flags & T139;
  assign T139 = ~ T140;
  assign T140 = 1'h1 << T165;
  assign T141 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T142;
  assign T142 = T51 ? T143 : 1'h0;
  assign T143 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T144;
  assign T144 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T145;
  assign T145 = 3'h5;
  assign io_inner_grant_bits_payload_client_xact_id = T146;
  assign T146 = xact_client_xact_id;
  assign T147 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T148;
  assign T148 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T168;
  assign T168 = {1'h0, init_client_id};
  assign T169 = T170[1'h0:1'h0];
  assign T170 = reset ? 2'h0 : T149;
  assign T149 = T21 ? io_inner_acquire_bits_header_src : T171;
  assign T171 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T150;
  assign T150 = T151 ? 1'h1 : T84;
  assign T151 = T88 & T152;
  assign T152 = io_outer_grant_valid & T153;
  assign T153 = T172 == 3'h5;
  assign T172 = {1'h0, io_outer_grant_bits_payload_client_xact_id};
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T81;
    end else if(T79) begin
      state <= T78;
    end else if(T76) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T155;
    init_sharer_cnt <= T161;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T141) begin
      probe_flags <= T138;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T169;
  end
endmodule

module AcquireTracker_5(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T154;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T155;
  wire[1:0] T156;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T157;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T158;
  wire T38;
  wire[1:0] T159;
  wire T39;
  wire[1:0] T160;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[3:0] T72;
  wire T73;
  reg  init_sharer_cnt;
  wire T161;
  wire[1:0] T162;
  wire[1:0] T74;
  wire[1:0] T163;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire[2:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg [25:0] xact_addr;
  wire[25:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T97;
  wire[2:0] T98;
  wire[2:0] T99;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T100;
  wire[5:0] T101;
  wire[5:0] T102;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T103;
  wire[2:0] T104;
  wire[2:0] T105;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T106;
  wire[511:0] T107;
  wire[511:0] T108;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T113;
  wire[25:0] T114;
  wire[25:0] T115;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T116;
  wire T117;
  wire T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[25:0] T135;
  wire[1:0] T164;
  wire T165;
  wire T166;
  reg [1:0] probe_flags;
  wire[1:0] T167;
  wire[1:0] T136;
  wire[1:0] T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire[3:0] T144;
  wire[2:0] T145;
  wire[1:0] T146;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T147;
  wire[511:0] T148;
  wire[1:0] T168;
  reg  init_client_id;
  wire T169;
  wire[1:0] T170;
  wire[1:0] T149;
  wire[1:0] T171;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire[2:0] T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T154 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T81 : T4;
  assign T4 = T79 ? T78 : T5;
  assign T5 = T76 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T155 = T156[1'h0:1'h0];
  assign T156 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T160 : T33;
  assign T33 = T52 ? T159 : T34;
  assign T34 = T21 ? T35 : T157;
  assign T157 = {1'h0, release_count};
  assign T35 = T158 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T158 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T159 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T160 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T75 ? T72 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = T73 ? 4'h1 : 4'h2;
  assign T73 = 1'h0 < init_sharer_cnt;
  assign T161 = T162[1'h0:1'h0];
  assign T162 = reset ? 2'h0 : T74;
  assign T74 = T21 ? 2'h2 : T163;
  assign T163 = {1'h0, init_sharer_cnt};
  assign T75 = xact_a_type == 3'h0;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h2 == state;
  assign T78 = pending_outer_read ? 3'h2 : 3'h4;
  assign T79 = T80 & io_outer_acquire_ready;
  assign T80 = 3'h3 == state;
  assign T81 = T82 ? 3'h5 : 3'h0;
  assign T82 = grant_type != 4'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_master_xact_id == 3'h6;
  assign T88 = 3'h5 == state;
  assign T89 = xact_addr == io_inner_release_bits_payload_addr;
  assign T90 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T91;
  assign T91 = T93 & T92;
  assign T92 = state != 3'h0;
  assign T93 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T94;
  assign T94 = T80 ? outer_write_acq_atomic_opcode : T95;
  assign T95 = T77 ? outer_read_atomic_opcode : T96;
  assign T96 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T97;
  assign T97 = T80 ? outer_write_acq_subword_addr : T98;
  assign T98 = T77 ? outer_read_subword_addr : T99;
  assign T99 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T100;
  assign T100 = T80 ? outer_write_acq_write_mask : T101;
  assign T101 = T77 ? outer_read_write_mask : T102;
  assign T102 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T103;
  assign T103 = T80 ? outer_write_acq_a_type : T104;
  assign T104 = T77 ? outer_read_a_type : T105;
  assign T105 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T106;
  assign T106 = T80 ? outer_write_acq_data : T107;
  assign T107 = T77 ? outer_read_data : T108;
  assign T108 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T109 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T110;
  assign T110 = T80 ? outer_write_acq_client_xact_id : T111;
  assign T111 = T77 ? outer_read_client_xact_id : T112;
  assign T112 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 2'h2;
  assign outer_read_client_xact_id = 2'h2;
  assign outer_write_acq_client_xact_id = 2'h2;
  assign io_outer_acquire_bits_payload_addr = T113;
  assign T113 = T80 ? outer_write_acq_addr : T114;
  assign T114 = T77 ? outer_read_addr : T115;
  assign T115 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T116;
  assign T116 = T80 ? 1'h1 : T117;
  assign T117 = T77 ? 1'h1 : T53;
  assign io_inner_release_ready = T118;
  assign T118 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T119;
  assign T119 = T120;
  assign T120 = T133 ? 2'h1 : T121;
  assign T121 = T132 ? 2'h0 : T122;
  assign T122 = T131 ? 2'h2 : T123;
  assign T123 = T130 ? 2'h0 : T124;
  assign T124 = T129 ? 2'h2 : T125;
  assign T125 = T128 ? 2'h0 : T126;
  assign T126 = T127 ? 2'h0 : 2'h2;
  assign T127 = xact_a_type == 3'h6;
  assign T128 = xact_a_type == 3'h5;
  assign T129 = xact_a_type == 3'h4;
  assign T130 = xact_a_type == 3'h3;
  assign T131 = xact_a_type == 3'h2;
  assign T132 = xact_a_type == 3'h1;
  assign T133 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T134;
  assign T134 = 3'h6;
  assign io_inner_probe_bits_payload_addr = T135;
  assign T135 = xact_addr;
  assign io_inner_probe_bits_header_dst = T164;
  assign T164 = {1'h0, T165};
  assign T165 = T166 == 1'h0;
  assign T166 = probe_flags[1'h0:1'h0];
  assign T167 = reset ? 2'h0 : T136;
  assign T136 = T141 ? T138 : T137;
  assign T137 = T21 ? probe_initial_flags : probe_flags;
  assign T138 = probe_flags & T139;
  assign T139 = ~ T140;
  assign T140 = 1'h1 << T165;
  assign T141 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T142;
  assign T142 = T51 ? T143 : 1'h0;
  assign T143 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T144;
  assign T144 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T145;
  assign T145 = 3'h6;
  assign io_inner_grant_bits_payload_client_xact_id = T146;
  assign T146 = xact_client_xact_id;
  assign T147 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T148;
  assign T148 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T168;
  assign T168 = {1'h0, init_client_id};
  assign T169 = T170[1'h0:1'h0];
  assign T170 = reset ? 2'h0 : T149;
  assign T149 = T21 ? io_inner_acquire_bits_header_src : T171;
  assign T171 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T150;
  assign T150 = T151 ? 1'h1 : T84;
  assign T151 = T88 & T152;
  assign T152 = io_outer_grant_valid & T153;
  assign T153 = T172 == 3'h6;
  assign T172 = {1'h0, io_outer_grant_bits_payload_client_xact_id};
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T81;
    end else if(T79) begin
      state <= T78;
    end else if(T76) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T155;
    init_sharer_cnt <= T161;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T141) begin
      probe_flags <= T138;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T169;
  end
endmodule

module AcquireTracker_6(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T154;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] probe_initial_flags;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire pending_outer_read;
  reg [2:0] xact_a_type;
  wire[2:0] T25;
  wire pending_outer_write;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg  release_count;
  wire T155;
  wire[1:0] T156;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T157;
  wire[1:0] T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T158;
  wire T38;
  wire[1:0] T159;
  wire T39;
  wire[1:0] T160;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire[3:0] grant_type;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[3:0] T72;
  wire T73;
  reg  init_sharer_cnt;
  wire T161;
  wire[1:0] T162;
  wire[1:0] T74;
  wire[1:0] T163;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire T79;
  wire T80;
  wire[2:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg [25:0] xact_addr;
  wire[25:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T97;
  wire[2:0] T98;
  wire[2:0] T99;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T100;
  wire[5:0] T101;
  wire[5:0] T102;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T103;
  wire[2:0] T104;
  wire[2:0] T105;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T106;
  wire[511:0] T107;
  wire[511:0] T108;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T113;
  wire[25:0] T114;
  wire[25:0] T115;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_acq_addr;
  wire T116;
  wire T117;
  wire T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] T124;
  wire[1:0] T125;
  wire[1:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[25:0] T135;
  wire[1:0] T164;
  wire T165;
  wire T166;
  reg [1:0] probe_flags;
  wire[1:0] T167;
  wire[1:0] T136;
  wire[1:0] T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire[3:0] T144;
  wire[2:0] T145;
  wire[1:0] T146;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T147;
  wire[511:0] T148;
  wire[1:0] T168;
  reg  init_client_id;
  wire T169;
  wire[1:0] T170;
  wire[1:0] T149;
  wire[1:0] T171;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire[2:0] T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T89 & T1;
  assign T1 = state != 3'h0;
  assign T154 = reset ? 3'h0 : T2;
  assign T2 = T85 ? 3'h0 : T3;
  assign T3 = T83 ? T81 : T4;
  assign T4 = T79 ? T78 : T5;
  assign T5 = T76 ? T58 : T6;
  assign T6 = T56 ? T54 : T7;
  assign T7 = T30 ? T23 : T8;
  assign T8 = T21 ? T9 : state;
  assign T9 = T18 ? 3'h1 : T10;
  assign T10 = T13 ? 3'h3 : T11;
  assign T11 = T12 ? 3'h2 : 3'h4;
  assign T12 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T13 = T15 | T14;
  assign T14 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T15 = T17 | T16;
  assign T16 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T17 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T18 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T19;
  assign T19 = ~ T20;
  assign T20 = io_tile_incoherent | 2'h0;
  assign T21 = T22 & io_inner_acquire_valid;
  assign T22 = 3'h0 == state;
  assign T23 = pending_outer_write ? 3'h3 : T24;
  assign T24 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = xact_a_type != 3'h3;
  assign T25 = T21 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T27 | T26;
  assign T26 = 3'h6 == xact_a_type;
  assign T27 = T29 | T28;
  assign T28 = 3'h5 == xact_a_type;
  assign T29 = 3'h3 == xact_a_type;
  assign T30 = T52 & T31;
  assign T31 = release_count == 1'h1;
  assign T155 = T156[1'h0:1'h0];
  assign T156 = reset ? 2'h0 : T32;
  assign T32 = T41 ? T160 : T33;
  assign T33 = T52 ? T159 : T34;
  assign T34 = T21 ? T35 : T157;
  assign T157 = {1'h0, release_count};
  assign T35 = T158 + T36;
  assign T36 = {1'h0, T37};
  assign T37 = probe_initial_flags[1'h1:1'h1];
  assign T158 = {1'h0, T38};
  assign T38 = probe_initial_flags[1'h0:1'h0];
  assign T159 = {1'h0, T39};
  assign T39 = release_count - 1'h1;
  assign T160 = {1'h0, T40};
  assign T40 = release_count - 1'h1;
  assign T41 = T50 & T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T45 | T44;
  assign T44 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T45 = T47 | T46;
  assign T46 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T47 = T49 | T48;
  assign T48 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T49 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T50 = T51 & io_inner_release_valid;
  assign T51 = 3'h1 == state;
  assign T52 = T53 & io_outer_acquire_ready;
  assign T53 = T50 & T43;
  assign T54 = pending_outer_write ? 3'h3 : T55;
  assign T55 = pending_outer_read ? 3'h2 : 3'h4;
  assign T56 = T41 & T57;
  assign T57 = release_count == 1'h1;
  assign T58 = T59 ? 3'h5 : 3'h0;
  assign T59 = grant_type != 4'h0;
  assign grant_type = T75 ? T72 : T60;
  assign T60 = T71 ? 4'h2 : T61;
  assign T61 = T70 ? 4'h3 : T62;
  assign T62 = T69 ? 4'h4 : T63;
  assign T63 = T68 ? 4'h6 : T64;
  assign T64 = T67 ? 4'h7 : T65;
  assign T65 = T66 ? 4'h8 : 4'h3;
  assign T66 = xact_a_type == 3'h6;
  assign T67 = xact_a_type == 3'h5;
  assign T68 = xact_a_type == 3'h4;
  assign T69 = xact_a_type == 3'h3;
  assign T70 = xact_a_type == 3'h2;
  assign T71 = xact_a_type == 3'h1;
  assign T72 = T73 ? 4'h1 : 4'h2;
  assign T73 = 1'h0 < init_sharer_cnt;
  assign T161 = T162[1'h0:1'h0];
  assign T162 = reset ? 2'h0 : T74;
  assign T74 = T21 ? 2'h2 : T163;
  assign T163 = {1'h0, init_sharer_cnt};
  assign T75 = xact_a_type == 3'h0;
  assign T76 = T77 & io_outer_acquire_ready;
  assign T77 = 3'h2 == state;
  assign T78 = pending_outer_read ? 3'h2 : 3'h4;
  assign T79 = T80 & io_outer_acquire_ready;
  assign T80 = 3'h3 == state;
  assign T81 = T82 ? 3'h5 : 3'h0;
  assign T82 = grant_type != 4'h0;
  assign T83 = T84 & io_inner_grant_ready;
  assign T84 = 3'h4 == state;
  assign T85 = T88 & T86;
  assign T86 = io_inner_finish_valid & T87;
  assign T87 = io_inner_finish_bits_payload_master_xact_id == 3'h7;
  assign T88 = 3'h5 == state;
  assign T89 = xact_addr == io_inner_release_bits_payload_addr;
  assign T90 = T21 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T91;
  assign T91 = T93 & T92;
  assign T92 = state != 3'h0;
  assign T93 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T94;
  assign T94 = T80 ? outer_write_acq_atomic_opcode : T95;
  assign T95 = T77 ? outer_read_atomic_opcode : T96;
  assign T96 = T53 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T97;
  assign T97 = T80 ? outer_write_acq_subword_addr : T98;
  assign T98 = T77 ? outer_read_subword_addr : T99;
  assign T99 = T53 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T100;
  assign T100 = T80 ? outer_write_acq_write_mask : T101;
  assign T101 = T77 ? outer_read_write_mask : T102;
  assign T102 = T53 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T103;
  assign T103 = T80 ? outer_write_acq_a_type : T104;
  assign T104 = T77 ? outer_read_a_type : T105;
  assign T105 = T53 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_read_a_type = 3'h2;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T106;
  assign T106 = T80 ? outer_write_acq_data : T107;
  assign T107 = T77 ? outer_read_data : T108;
  assign T108 = T53 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_read_data = 512'h0;
  assign outer_write_acq_data = xact_data;
  assign T109 = T21 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T110;
  assign T110 = T80 ? outer_write_acq_client_xact_id : T111;
  assign T111 = T77 ? outer_read_client_xact_id : T112;
  assign T112 = T53 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 2'h3;
  assign outer_read_client_xact_id = 2'h3;
  assign outer_write_acq_client_xact_id = 2'h3;
  assign io_outer_acquire_bits_payload_addr = T113;
  assign T113 = T80 ? outer_write_acq_addr : T114;
  assign T114 = T77 ? outer_read_addr : T115;
  assign T115 = T53 ? outer_write_rel_addr : outer_read_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T116;
  assign T116 = T80 ? 1'h1 : T117;
  assign T117 = T77 ? 1'h1 : T53;
  assign io_inner_release_ready = T118;
  assign T118 = T41 ? 1'h1 : T52;
  assign io_inner_probe_bits_payload_p_type = T119;
  assign T119 = T120;
  assign T120 = T133 ? 2'h1 : T121;
  assign T121 = T132 ? 2'h0 : T122;
  assign T122 = T131 ? 2'h2 : T123;
  assign T123 = T130 ? 2'h0 : T124;
  assign T124 = T129 ? 2'h2 : T125;
  assign T125 = T128 ? 2'h0 : T126;
  assign T126 = T127 ? 2'h0 : 2'h2;
  assign T127 = xact_a_type == 3'h6;
  assign T128 = xact_a_type == 3'h5;
  assign T129 = xact_a_type == 3'h4;
  assign T130 = xact_a_type == 3'h3;
  assign T131 = xact_a_type == 3'h2;
  assign T132 = xact_a_type == 3'h1;
  assign T133 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T134;
  assign T134 = 3'h7;
  assign io_inner_probe_bits_payload_addr = T135;
  assign T135 = xact_addr;
  assign io_inner_probe_bits_header_dst = T164;
  assign T164 = {1'h0, T165};
  assign T165 = T166 == 1'h0;
  assign T166 = probe_flags[1'h0:1'h0];
  assign T167 = reset ? 2'h0 : T136;
  assign T136 = T141 ? T138 : T137;
  assign T137 = T21 ? probe_initial_flags : probe_flags;
  assign T138 = probe_flags & T139;
  assign T139 = ~ T140;
  assign T140 = 1'h1 << T165;
  assign T141 = T51 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T142;
  assign T142 = T51 ? T143 : 1'h0;
  assign T143 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T144;
  assign T144 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T145;
  assign T145 = 3'h7;
  assign io_inner_grant_bits_payload_client_xact_id = T146;
  assign T146 = xact_client_xact_id;
  assign T147 = T21 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T148;
  assign T148 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T168;
  assign T168 = {1'h0, init_client_id};
  assign T169 = T170[1'h0:1'h0];
  assign T170 = reset ? 2'h0 : T149;
  assign T149 = T21 ? io_inner_acquire_bits_header_src : T171;
  assign T171 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T150;
  assign T150 = T151 ? 1'h1 : T84;
  assign T151 = T88 & T152;
  assign T152 = io_outer_grant_valid & T153;
  assign T153 = T172 == 3'h7;
  assign T172 = {1'h0, io_outer_grant_bits_payload_client_xact_id};
  assign io_inner_acquire_ready = T22;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T85) begin
      state <= 3'h0;
    end else if(T83) begin
      state <= T81;
    end else if(T79) begin
      state <= T78;
    end else if(T76) begin
      state <= T58;
    end else if(T56) begin
      state <= T54;
    end else if(T30) begin
      state <= T23;
    end else if(T21) begin
      state <= T9;
    end
    if(T21) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T155;
    init_sharer_cnt <= T161;
    if(T21) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T21) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T141) begin
      probe_flags <= T138;
    end else if(T21) begin
      probe_flags <= probe_initial_flags;
    end
    if(T21) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T169;
  end
endmodule

module Arbiter_11(
    output io_in_7_ready,
    input  io_in_7_valid,
    input  io_in_7_bits,
    output io_in_6_ready,
    input  io_in_6_valid,
    input  io_in_6_bits,
    output io_in_5_ready,
    input  io_in_5_valid,
    input  io_in_5_bits,
    output io_in_4_ready,
    input  io_in_4_valid,
    input  io_in_4_bits,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits : io_in_0_bits;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits : io_in_2_bits;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits : io_in_4_bits;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits : io_in_6_bits;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_valid = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_valid : io_in_0_valid;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_valid : io_in_2_valid;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_valid : io_in_4_valid;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_valid : io_in_6_valid;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T37;
  assign T37 = T38 & io_out_ready;
  assign T38 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T41 ^ 1'h1;
  assign T41 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T42;
  assign T42 = T43 & io_out_ready;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T45 | io_in_2_valid;
  assign T45 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T46;
  assign T46 = T47 & io_out_ready;
  assign T47 = T48 ^ 1'h1;
  assign T48 = T49 | io_in_3_valid;
  assign T49 = T50 | io_in_2_valid;
  assign T50 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T54 | io_in_4_valid;
  assign T54 = T55 | io_in_3_valid;
  assign T55 = T56 | io_in_2_valid;
  assign T56 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T57;
  assign T57 = T58 & io_out_ready;
  assign T58 = T59 ^ 1'h1;
  assign T59 = T60 | io_in_5_valid;
  assign T60 = T61 | io_in_4_valid;
  assign T61 = T62 | io_in_3_valid;
  assign T62 = T63 | io_in_2_valid;
  assign T63 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_6_valid;
  assign T67 = T68 | io_in_5_valid;
  assign T68 = T69 | io_in_4_valid;
  assign T69 = T70 | io_in_3_valid;
  assign T70 = T71 | io_in_2_valid;
  assign T71 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_12(
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [2:0] io_in_7_bits_payload_master_xact_id,
    input [1:0] io_in_7_bits_payload_p_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [2:0] io_in_6_bits_payload_master_xact_id,
    input [1:0] io_in_6_bits_payload_p_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [2:0] io_in_5_bits_payload_master_xact_id,
    input [1:0] io_in_5_bits_payload_p_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [2:0] io_in_4_bits_payload_master_xact_id,
    input [1:0] io_in_4_bits_payload_p_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [2:0] io_in_3_bits_payload_master_xact_id,
    input [1:0] io_in_3_bits_payload_p_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_out_bits_payload_p_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire[2:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire[25:0] T37;
  wire[25:0] T38;
  wire[25:0] T39;
  wire T40;
  wire[25:0] T41;
  wire T42;
  wire T43;
  wire[25:0] T44;
  wire[25:0] T45;
  wire T46;
  wire[25:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[1:0] T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits_payload_p_type = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits_payload_p_type : io_in_2_bits_payload_p_type;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits_payload_p_type : io_in_4_bits_payload_p_type;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits_payload_p_type : io_in_6_bits_payload_p_type;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_bits_payload_master_xact_id = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_out_bits_payload_addr = T37;
  assign T37 = T50 ? T44 : T38;
  assign T38 = T43 ? T41 : T39;
  assign T39 = T40 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T40 = T12[1'h0:1'h0];
  assign T41 = T42 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T42 = T12[1'h0:1'h0];
  assign T43 = T12[1'h1:1'h1];
  assign T44 = T49 ? T47 : T45;
  assign T45 = T46 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T46 = T12[1'h0:1'h0];
  assign T47 = T48 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T48 = T12[1'h0:1'h0];
  assign T49 = T12[1'h1:1'h1];
  assign T50 = T12[2'h2:2'h2];
  assign io_out_bits_header_dst = T51;
  assign T51 = T64 ? T58 : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T54 = T12[1'h0:1'h0];
  assign T55 = T56 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T56 = T12[1'h0:1'h0];
  assign T57 = T12[1'h1:1'h1];
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T60 = T12[1'h0:1'h0];
  assign T61 = T62 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T62 = T12[1'h0:1'h0];
  assign T63 = T12[1'h1:1'h1];
  assign T64 = T12[2'h2:2'h2];
  assign io_out_bits_header_src = T65;
  assign T65 = T78 ? T72 : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T68 = T12[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T70 = T12[1'h0:1'h0];
  assign T71 = T12[1'h1:1'h1];
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T74 = T12[1'h0:1'h0];
  assign T75 = T76 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T76 = T12[1'h0:1'h0];
  assign T77 = T12[1'h1:1'h1];
  assign T78 = T12[2'h2:2'h2];
  assign io_out_valid = T79;
  assign T79 = T92 ? T86 : T80;
  assign T80 = T85 ? T83 : T81;
  assign T81 = T82 ? io_in_1_valid : io_in_0_valid;
  assign T82 = T12[1'h0:1'h0];
  assign T83 = T84 ? io_in_3_valid : io_in_2_valid;
  assign T84 = T12[1'h0:1'h0];
  assign T85 = T12[1'h1:1'h1];
  assign T86 = T91 ? T89 : T87;
  assign T87 = T88 ? io_in_5_valid : io_in_4_valid;
  assign T88 = T12[1'h0:1'h0];
  assign T89 = T90 ? io_in_7_valid : io_in_6_valid;
  assign T90 = T12[1'h0:1'h0];
  assign T91 = T12[1'h1:1'h1];
  assign T92 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T93;
  assign T93 = T94 & io_out_ready;
  assign T94 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T95;
  assign T95 = T96 & io_out_ready;
  assign T96 = T97 ^ 1'h1;
  assign T97 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T98;
  assign T98 = T99 & io_out_ready;
  assign T99 = T100 ^ 1'h1;
  assign T100 = T101 | io_in_2_valid;
  assign T101 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T102;
  assign T102 = T103 & io_out_ready;
  assign T103 = T104 ^ 1'h1;
  assign T104 = T105 | io_in_3_valid;
  assign T105 = T106 | io_in_2_valid;
  assign T106 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T107;
  assign T107 = T108 & io_out_ready;
  assign T108 = T109 ^ 1'h1;
  assign T109 = T110 | io_in_4_valid;
  assign T110 = T111 | io_in_3_valid;
  assign T111 = T112 | io_in_2_valid;
  assign T112 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T113;
  assign T113 = T114 & io_out_ready;
  assign T114 = T115 ^ 1'h1;
  assign T115 = T116 | io_in_5_valid;
  assign T116 = T117 | io_in_4_valid;
  assign T117 = T118 | io_in_3_valid;
  assign T118 = T119 | io_in_2_valid;
  assign T119 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T120;
  assign T120 = T121 & io_out_ready;
  assign T121 = T122 ^ 1'h1;
  assign T122 = T123 | io_in_6_valid;
  assign T123 = T124 | io_in_5_valid;
  assign T124 = T125 | io_in_4_valid;
  assign T125 = T126 | io_in_3_valid;
  assign T126 = T127 | io_in_2_valid;
  assign T127 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_13(
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [511:0] io_in_7_bits_payload_data,
    input [1:0] io_in_7_bits_payload_client_xact_id,
    input [2:0] io_in_7_bits_payload_master_xact_id,
    input [3:0] io_in_7_bits_payload_g_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [511:0] io_in_6_bits_payload_data,
    input [1:0] io_in_6_bits_payload_client_xact_id,
    input [2:0] io_in_6_bits_payload_master_xact_id,
    input [3:0] io_in_6_bits_payload_g_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [511:0] io_in_5_bits_payload_data,
    input [1:0] io_in_5_bits_payload_client_xact_id,
    input [2:0] io_in_5_bits_payload_master_xact_id,
    input [3:0] io_in_5_bits_payload_g_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [511:0] io_in_4_bits_payload_data,
    input [1:0] io_in_4_bits_payload_client_xact_id,
    input [2:0] io_in_4_bits_payload_master_xact_id,
    input [3:0] io_in_4_bits_payload_g_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [511:0] io_in_3_bits_payload_data,
    input [1:0] io_in_3_bits_payload_client_xact_id,
    input [2:0] io_in_3_bits_payload_master_xact_id,
    input [3:0] io_in_3_bits_payload_g_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire T11;
  wire[2:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire T18;
  wire[3:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[511:0] T51;
  wire[511:0] T52;
  wire[511:0] T53;
  wire T54;
  wire[511:0] T55;
  wire T56;
  wire T57;
  wire[511:0] T58;
  wire[511:0] T59;
  wire T60;
  wire[511:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[1:0] T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire[1:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits_payload_g_type = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits_payload_g_type : io_in_2_bits_payload_g_type;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits_payload_g_type : io_in_4_bits_payload_g_type;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits_payload_g_type : io_in_6_bits_payload_g_type;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_bits_payload_master_xact_id = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T37;
  assign T37 = T50 ? T44 : T38;
  assign T38 = T43 ? T41 : T39;
  assign T39 = T40 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T40 = T12[1'h0:1'h0];
  assign T41 = T42 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T42 = T12[1'h0:1'h0];
  assign T43 = T12[1'h1:1'h1];
  assign T44 = T49 ? T47 : T45;
  assign T45 = T46 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T46 = T12[1'h0:1'h0];
  assign T47 = T48 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T48 = T12[1'h0:1'h0];
  assign T49 = T12[1'h1:1'h1];
  assign T50 = T12[2'h2:2'h2];
  assign io_out_bits_payload_data = T51;
  assign T51 = T64 ? T58 : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T54 = T12[1'h0:1'h0];
  assign T55 = T56 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T56 = T12[1'h0:1'h0];
  assign T57 = T12[1'h1:1'h1];
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T60 = T12[1'h0:1'h0];
  assign T61 = T62 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T62 = T12[1'h0:1'h0];
  assign T63 = T12[1'h1:1'h1];
  assign T64 = T12[2'h2:2'h2];
  assign io_out_bits_header_dst = T65;
  assign T65 = T78 ? T72 : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T68 = T12[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T70 = T12[1'h0:1'h0];
  assign T71 = T12[1'h1:1'h1];
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T74 = T12[1'h0:1'h0];
  assign T75 = T76 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T76 = T12[1'h0:1'h0];
  assign T77 = T12[1'h1:1'h1];
  assign T78 = T12[2'h2:2'h2];
  assign io_out_bits_header_src = T79;
  assign T79 = T92 ? T86 : T80;
  assign T80 = T85 ? T83 : T81;
  assign T81 = T82 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T82 = T12[1'h0:1'h0];
  assign T83 = T84 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T84 = T12[1'h0:1'h0];
  assign T85 = T12[1'h1:1'h1];
  assign T86 = T91 ? T89 : T87;
  assign T87 = T88 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T88 = T12[1'h0:1'h0];
  assign T89 = T90 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T90 = T12[1'h0:1'h0];
  assign T91 = T12[1'h1:1'h1];
  assign T92 = T12[2'h2:2'h2];
  assign io_out_valid = T93;
  assign T93 = T106 ? T100 : T94;
  assign T94 = T99 ? T97 : T95;
  assign T95 = T96 ? io_in_1_valid : io_in_0_valid;
  assign T96 = T12[1'h0:1'h0];
  assign T97 = T98 ? io_in_3_valid : io_in_2_valid;
  assign T98 = T12[1'h0:1'h0];
  assign T99 = T12[1'h1:1'h1];
  assign T100 = T105 ? T103 : T101;
  assign T101 = T102 ? io_in_5_valid : io_in_4_valid;
  assign T102 = T12[1'h0:1'h0];
  assign T103 = T104 ? io_in_7_valid : io_in_6_valid;
  assign T104 = T12[1'h0:1'h0];
  assign T105 = T12[1'h1:1'h1];
  assign T106 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T107;
  assign T107 = T108 & io_out_ready;
  assign T108 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T109;
  assign T109 = T110 & io_out_ready;
  assign T110 = T111 ^ 1'h1;
  assign T111 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T112;
  assign T112 = T113 & io_out_ready;
  assign T113 = T114 ^ 1'h1;
  assign T114 = T115 | io_in_2_valid;
  assign T115 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T116;
  assign T116 = T117 & io_out_ready;
  assign T117 = T118 ^ 1'h1;
  assign T118 = T119 | io_in_3_valid;
  assign T119 = T120 | io_in_2_valid;
  assign T120 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T121;
  assign T121 = T122 & io_out_ready;
  assign T122 = T123 ^ 1'h1;
  assign T123 = T124 | io_in_4_valid;
  assign T124 = T125 | io_in_3_valid;
  assign T125 = T126 | io_in_2_valid;
  assign T126 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T127;
  assign T127 = T128 & io_out_ready;
  assign T128 = T129 ^ 1'h1;
  assign T129 = T130 | io_in_5_valid;
  assign T130 = T131 | io_in_4_valid;
  assign T131 = T132 | io_in_3_valid;
  assign T132 = T133 | io_in_2_valid;
  assign T133 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T134;
  assign T134 = T135 & io_out_ready;
  assign T135 = T136 ^ 1'h1;
  assign T136 = T137 | io_in_6_valid;
  assign T137 = T138 | io_in_5_valid;
  assign T138 = T139 | io_in_4_valid;
  assign T139 = T140 | io_in_3_valid;
  assign T140 = T141 | io_in_2_valid;
  assign T141 = io_in_0_valid | io_in_1_valid;
endmodule

module RRArbiter_3(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [1:0] io_in_7_bits_payload_client_xact_id,
    input [511:0] io_in_7_bits_payload_data,
    input [2:0] io_in_7_bits_payload_a_type,
    input [5:0] io_in_7_bits_payload_write_mask,
    input [2:0] io_in_7_bits_payload_subword_addr,
    input [3:0] io_in_7_bits_payload_atomic_opcode,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [1:0] io_in_6_bits_payload_client_xact_id,
    input [511:0] io_in_6_bits_payload_data,
    input [2:0] io_in_6_bits_payload_a_type,
    input [5:0] io_in_6_bits_payload_write_mask,
    input [2:0] io_in_6_bits_payload_subword_addr,
    input [3:0] io_in_6_bits_payload_atomic_opcode,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [1:0] io_in_5_bits_payload_client_xact_id,
    input [511:0] io_in_5_bits_payload_data,
    input [2:0] io_in_5_bits_payload_a_type,
    input [5:0] io_in_5_bits_payload_write_mask,
    input [2:0] io_in_5_bits_payload_subword_addr,
    input [3:0] io_in_5_bits_payload_atomic_opcode,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [1:0] io_in_4_bits_payload_client_xact_id,
    input [511:0] io_in_4_bits_payload_data,
    input [2:0] io_in_4_bits_payload_a_type,
    input [5:0] io_in_4_bits_payload_write_mask,
    input [2:0] io_in_4_bits_payload_subword_addr,
    input [3:0] io_in_4_bits_payload_atomic_opcode,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [1:0] io_in_3_bits_payload_client_xact_id,
    input [511:0] io_in_3_bits_payload_data,
    input [2:0] io_in_3_bits_payload_a_type,
    input [5:0] io_in_3_bits_payload_write_mask,
    input [2:0] io_in_3_bits_payload_subword_addr,
    input [3:0] io_in_3_bits_payload_atomic_opcode,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  reg [2:0] R17;
  wire[2:0] T340;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire T35;
  wire[2:0] T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire[3:0] T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire[2:0] T47;
  wire[2:0] T48;
  wire[2:0] T49;
  wire T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;
  wire[2:0] T55;
  wire T56;
  wire[2:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[5:0] T61;
  wire[5:0] T62;
  wire[5:0] T63;
  wire T64;
  wire[5:0] T65;
  wire T66;
  wire T67;
  wire[5:0] T68;
  wire[5:0] T69;
  wire T70;
  wire[5:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire[2:0] T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire T78;
  wire[2:0] T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire[2:0] T83;
  wire T84;
  wire[2:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[511:0] T89;
  wire[511:0] T90;
  wire[511:0] T91;
  wire T92;
  wire[511:0] T93;
  wire T94;
  wire T95;
  wire[511:0] T96;
  wire[511:0] T97;
  wire T98;
  wire[511:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  wire[1:0] T107;
  wire T108;
  wire T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire T112;
  wire[1:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[25:0] T117;
  wire[25:0] T118;
  wire[25:0] T119;
  wire T120;
  wire[25:0] T121;
  wire T122;
  wire T123;
  wire[25:0] T124;
  wire[25:0] T125;
  wire T126;
  wire[25:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire[1:0] T138;
  wire[1:0] T139;
  wire T140;
  wire[1:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[1:0] T145;
  wire[1:0] T146;
  wire[1:0] T147;
  wire T148;
  wire[1:0] T149;
  wire T150;
  wire T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T30 ? 3'h1 : T2;
  assign T2 = T28 ? 3'h2 : T3;
  assign T3 = T26 ? 3'h3 : T4;
  assign T4 = T24 ? 3'h4 : T5;
  assign T5 = T22 ? 3'h5 : T6;
  assign T6 = T20 ? 3'h6 : T7;
  assign T7 = T15 ? 3'h7 : T8;
  assign T8 = io_in_0_valid ? 3'h0 : T9;
  assign T9 = io_in_1_valid ? 3'h1 : T10;
  assign T10 = io_in_2_valid ? 3'h2 : T11;
  assign T11 = io_in_3_valid ? 3'h3 : T12;
  assign T12 = io_in_4_valid ? 3'h4 : T13;
  assign T13 = io_in_5_valid ? 3'h5 : T14;
  assign T14 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T15 = io_in_7_valid & T16;
  assign T16 = R17 < 3'h7;
  assign T340 = reset ? 3'h0 : T18;
  assign T18 = T19 ? T0 : R17;
  assign T19 = io_out_ready & io_out_valid;
  assign T20 = io_in_6_valid & T21;
  assign T21 = R17 < 3'h6;
  assign T22 = io_in_5_valid & T23;
  assign T23 = R17 < 3'h5;
  assign T24 = io_in_4_valid & T25;
  assign T25 = R17 < 3'h4;
  assign T26 = io_in_3_valid & T27;
  assign T27 = R17 < 3'h3;
  assign T28 = io_in_2_valid & T29;
  assign T29 = R17 < 3'h2;
  assign T30 = io_in_1_valid & T31;
  assign T31 = R17 < 3'h1;
  assign io_out_bits_payload_atomic_opcode = T32;
  assign T32 = T46 ? T40 : T33;
  assign T33 = T39 ? T37 : T34;
  assign T34 = T35 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T35 = T36[1'h0:1'h0];
  assign T36 = T0;
  assign T37 = T38 ? io_in_3_bits_payload_atomic_opcode : io_in_2_bits_payload_atomic_opcode;
  assign T38 = T36[1'h0:1'h0];
  assign T39 = T36[1'h1:1'h1];
  assign T40 = T45 ? T43 : T41;
  assign T41 = T42 ? io_in_5_bits_payload_atomic_opcode : io_in_4_bits_payload_atomic_opcode;
  assign T42 = T36[1'h0:1'h0];
  assign T43 = T44 ? io_in_7_bits_payload_atomic_opcode : io_in_6_bits_payload_atomic_opcode;
  assign T44 = T36[1'h0:1'h0];
  assign T45 = T36[1'h1:1'h1];
  assign T46 = T36[2'h2:2'h2];
  assign io_out_bits_payload_subword_addr = T47;
  assign T47 = T60 ? T54 : T48;
  assign T48 = T53 ? T51 : T49;
  assign T49 = T50 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign T50 = T36[1'h0:1'h0];
  assign T51 = T52 ? io_in_3_bits_payload_subword_addr : io_in_2_bits_payload_subword_addr;
  assign T52 = T36[1'h0:1'h0];
  assign T53 = T36[1'h1:1'h1];
  assign T54 = T59 ? T57 : T55;
  assign T55 = T56 ? io_in_5_bits_payload_subword_addr : io_in_4_bits_payload_subword_addr;
  assign T56 = T36[1'h0:1'h0];
  assign T57 = T58 ? io_in_7_bits_payload_subword_addr : io_in_6_bits_payload_subword_addr;
  assign T58 = T36[1'h0:1'h0];
  assign T59 = T36[1'h1:1'h1];
  assign T60 = T36[2'h2:2'h2];
  assign io_out_bits_payload_write_mask = T61;
  assign T61 = T74 ? T68 : T62;
  assign T62 = T67 ? T65 : T63;
  assign T63 = T64 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign T64 = T36[1'h0:1'h0];
  assign T65 = T66 ? io_in_3_bits_payload_write_mask : io_in_2_bits_payload_write_mask;
  assign T66 = T36[1'h0:1'h0];
  assign T67 = T36[1'h1:1'h1];
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_5_bits_payload_write_mask : io_in_4_bits_payload_write_mask;
  assign T70 = T36[1'h0:1'h0];
  assign T71 = T72 ? io_in_7_bits_payload_write_mask : io_in_6_bits_payload_write_mask;
  assign T72 = T36[1'h0:1'h0];
  assign T73 = T36[1'h1:1'h1];
  assign T74 = T36[2'h2:2'h2];
  assign io_out_bits_payload_a_type = T75;
  assign T75 = T88 ? T82 : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T78 = T36[1'h0:1'h0];
  assign T79 = T80 ? io_in_3_bits_payload_a_type : io_in_2_bits_payload_a_type;
  assign T80 = T36[1'h0:1'h0];
  assign T81 = T36[1'h1:1'h1];
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_5_bits_payload_a_type : io_in_4_bits_payload_a_type;
  assign T84 = T36[1'h0:1'h0];
  assign T85 = T86 ? io_in_7_bits_payload_a_type : io_in_6_bits_payload_a_type;
  assign T86 = T36[1'h0:1'h0];
  assign T87 = T36[1'h1:1'h1];
  assign T88 = T36[2'h2:2'h2];
  assign io_out_bits_payload_data = T89;
  assign T89 = T102 ? T96 : T90;
  assign T90 = T95 ? T93 : T91;
  assign T91 = T92 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T92 = T36[1'h0:1'h0];
  assign T93 = T94 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T94 = T36[1'h0:1'h0];
  assign T95 = T36[1'h1:1'h1];
  assign T96 = T101 ? T99 : T97;
  assign T97 = T98 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T98 = T36[1'h0:1'h0];
  assign T99 = T100 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T100 = T36[1'h0:1'h0];
  assign T101 = T36[1'h1:1'h1];
  assign T102 = T36[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T103;
  assign T103 = T116 ? T110 : T104;
  assign T104 = T109 ? T107 : T105;
  assign T105 = T106 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T106 = T36[1'h0:1'h0];
  assign T107 = T108 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T108 = T36[1'h0:1'h0];
  assign T109 = T36[1'h1:1'h1];
  assign T110 = T115 ? T113 : T111;
  assign T111 = T112 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T112 = T36[1'h0:1'h0];
  assign T113 = T114 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T114 = T36[1'h0:1'h0];
  assign T115 = T36[1'h1:1'h1];
  assign T116 = T36[2'h2:2'h2];
  assign io_out_bits_payload_addr = T117;
  assign T117 = T130 ? T124 : T118;
  assign T118 = T123 ? T121 : T119;
  assign T119 = T120 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T120 = T36[1'h0:1'h0];
  assign T121 = T122 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T122 = T36[1'h0:1'h0];
  assign T123 = T36[1'h1:1'h1];
  assign T124 = T129 ? T127 : T125;
  assign T125 = T126 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T126 = T36[1'h0:1'h0];
  assign T127 = T128 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T128 = T36[1'h0:1'h0];
  assign T129 = T36[1'h1:1'h1];
  assign T130 = T36[2'h2:2'h2];
  assign io_out_bits_header_dst = T131;
  assign T131 = T144 ? T138 : T132;
  assign T132 = T137 ? T135 : T133;
  assign T133 = T134 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T134 = T36[1'h0:1'h0];
  assign T135 = T136 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T136 = T36[1'h0:1'h0];
  assign T137 = T36[1'h1:1'h1];
  assign T138 = T143 ? T141 : T139;
  assign T139 = T140 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T140 = T36[1'h0:1'h0];
  assign T141 = T142 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T142 = T36[1'h0:1'h0];
  assign T143 = T36[1'h1:1'h1];
  assign T144 = T36[2'h2:2'h2];
  assign io_out_bits_header_src = T145;
  assign T145 = T158 ? T152 : T146;
  assign T146 = T151 ? T149 : T147;
  assign T147 = T148 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T148 = T36[1'h0:1'h0];
  assign T149 = T150 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T150 = T36[1'h0:1'h0];
  assign T151 = T36[1'h1:1'h1];
  assign T152 = T157 ? T155 : T153;
  assign T153 = T154 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T154 = T36[1'h0:1'h0];
  assign T155 = T156 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T156 = T36[1'h0:1'h0];
  assign T157 = T36[1'h1:1'h1];
  assign T158 = T36[2'h2:2'h2];
  assign io_out_valid = T159;
  assign T159 = T172 ? T166 : T160;
  assign T160 = T165 ? T163 : T161;
  assign T161 = T162 ? io_in_1_valid : io_in_0_valid;
  assign T162 = T36[1'h0:1'h0];
  assign T163 = T164 ? io_in_3_valid : io_in_2_valid;
  assign T164 = T36[1'h0:1'h0];
  assign T165 = T36[1'h1:1'h1];
  assign T166 = T171 ? T169 : T167;
  assign T167 = T168 ? io_in_5_valid : io_in_4_valid;
  assign T168 = T36[1'h0:1'h0];
  assign T169 = T170 ? io_in_7_valid : io_in_6_valid;
  assign T170 = T36[1'h0:1'h0];
  assign T171 = T36[1'h1:1'h1];
  assign T172 = T36[2'h2:2'h2];
  assign io_in_0_ready = T173;
  assign T173 = T174 & io_out_ready;
  assign T174 = T199 | T175;
  assign T175 = T176 ^ 1'h1;
  assign T176 = T179 | T177;
  assign T177 = io_in_7_valid & T178;
  assign T178 = R17 < 3'h7;
  assign T179 = T182 | T180;
  assign T180 = io_in_6_valid & T181;
  assign T181 = R17 < 3'h6;
  assign T182 = T185 | T183;
  assign T183 = io_in_5_valid & T184;
  assign T184 = R17 < 3'h5;
  assign T185 = T188 | T186;
  assign T186 = io_in_4_valid & T187;
  assign T187 = R17 < 3'h4;
  assign T188 = T191 | T189;
  assign T189 = io_in_3_valid & T190;
  assign T190 = R17 < 3'h3;
  assign T191 = T194 | T192;
  assign T192 = io_in_2_valid & T193;
  assign T193 = R17 < 3'h2;
  assign T194 = T197 | T195;
  assign T195 = io_in_1_valid & T196;
  assign T196 = R17 < 3'h1;
  assign T197 = io_in_0_valid & T198;
  assign T198 = R17 < 3'h0;
  assign T199 = R17 < 3'h0;
  assign io_in_1_ready = T200;
  assign T200 = T201 & io_out_ready;
  assign T201 = T211 | T202;
  assign T202 = T203 ^ 1'h1;
  assign T203 = T204 | io_in_0_valid;
  assign T204 = T205 | T177;
  assign T205 = T206 | T180;
  assign T206 = T207 | T183;
  assign T207 = T208 | T186;
  assign T208 = T209 | T189;
  assign T209 = T210 | T192;
  assign T210 = T197 | T195;
  assign T211 = T213 & T212;
  assign T212 = R17 < 3'h1;
  assign T213 = T197 ^ 1'h1;
  assign io_in_2_ready = T214;
  assign T214 = T215 & io_out_ready;
  assign T215 = T226 | T216;
  assign T216 = T217 ^ 1'h1;
  assign T217 = T218 | io_in_1_valid;
  assign T218 = T219 | io_in_0_valid;
  assign T219 = T220 | T177;
  assign T220 = T221 | T180;
  assign T221 = T222 | T183;
  assign T222 = T223 | T186;
  assign T223 = T224 | T189;
  assign T224 = T225 | T192;
  assign T225 = T197 | T195;
  assign T226 = T228 & T227;
  assign T227 = R17 < 3'h2;
  assign T228 = T229 ^ 1'h1;
  assign T229 = T197 | T195;
  assign io_in_3_ready = T230;
  assign T230 = T231 & io_out_ready;
  assign T231 = T243 | T232;
  assign T232 = T233 ^ 1'h1;
  assign T233 = T234 | io_in_2_valid;
  assign T234 = T235 | io_in_1_valid;
  assign T235 = T236 | io_in_0_valid;
  assign T236 = T237 | T177;
  assign T237 = T238 | T180;
  assign T238 = T239 | T183;
  assign T239 = T240 | T186;
  assign T240 = T241 | T189;
  assign T241 = T242 | T192;
  assign T242 = T197 | T195;
  assign T243 = T245 & T244;
  assign T244 = R17 < 3'h3;
  assign T245 = T246 ^ 1'h1;
  assign T246 = T247 | T192;
  assign T247 = T197 | T195;
  assign io_in_4_ready = T248;
  assign T248 = T249 & io_out_ready;
  assign T249 = T262 | T250;
  assign T250 = T251 ^ 1'h1;
  assign T251 = T252 | io_in_3_valid;
  assign T252 = T253 | io_in_2_valid;
  assign T253 = T254 | io_in_1_valid;
  assign T254 = T255 | io_in_0_valid;
  assign T255 = T256 | T177;
  assign T256 = T257 | T180;
  assign T257 = T258 | T183;
  assign T258 = T259 | T186;
  assign T259 = T260 | T189;
  assign T260 = T261 | T192;
  assign T261 = T197 | T195;
  assign T262 = T264 & T263;
  assign T263 = R17 < 3'h4;
  assign T264 = T265 ^ 1'h1;
  assign T265 = T266 | T189;
  assign T266 = T267 | T192;
  assign T267 = T197 | T195;
  assign io_in_5_ready = T268;
  assign T268 = T269 & io_out_ready;
  assign T269 = T283 | T270;
  assign T270 = T271 ^ 1'h1;
  assign T271 = T272 | io_in_4_valid;
  assign T272 = T273 | io_in_3_valid;
  assign T273 = T274 | io_in_2_valid;
  assign T274 = T275 | io_in_1_valid;
  assign T275 = T276 | io_in_0_valid;
  assign T276 = T277 | T177;
  assign T277 = T278 | T180;
  assign T278 = T279 | T183;
  assign T279 = T280 | T186;
  assign T280 = T281 | T189;
  assign T281 = T282 | T192;
  assign T282 = T197 | T195;
  assign T283 = T285 & T284;
  assign T284 = R17 < 3'h5;
  assign T285 = T286 ^ 1'h1;
  assign T286 = T287 | T186;
  assign T287 = T288 | T189;
  assign T288 = T289 | T192;
  assign T289 = T197 | T195;
  assign io_in_6_ready = T290;
  assign T290 = T291 & io_out_ready;
  assign T291 = T306 | T292;
  assign T292 = T293 ^ 1'h1;
  assign T293 = T294 | io_in_5_valid;
  assign T294 = T295 | io_in_4_valid;
  assign T295 = T296 | io_in_3_valid;
  assign T296 = T297 | io_in_2_valid;
  assign T297 = T298 | io_in_1_valid;
  assign T298 = T299 | io_in_0_valid;
  assign T299 = T300 | T177;
  assign T300 = T301 | T180;
  assign T301 = T302 | T183;
  assign T302 = T303 | T186;
  assign T303 = T304 | T189;
  assign T304 = T305 | T192;
  assign T305 = T197 | T195;
  assign T306 = T308 & T307;
  assign T307 = R17 < 3'h6;
  assign T308 = T309 ^ 1'h1;
  assign T309 = T310 | T183;
  assign T310 = T311 | T186;
  assign T311 = T312 | T189;
  assign T312 = T313 | T192;
  assign T313 = T197 | T195;
  assign io_in_7_ready = T314;
  assign T314 = T315 & io_out_ready;
  assign T315 = T331 | T316;
  assign T316 = T317 ^ 1'h1;
  assign T317 = T318 | io_in_6_valid;
  assign T318 = T319 | io_in_5_valid;
  assign T319 = T320 | io_in_4_valid;
  assign T320 = T321 | io_in_3_valid;
  assign T321 = T322 | io_in_2_valid;
  assign T322 = T323 | io_in_1_valid;
  assign T323 = T324 | io_in_0_valid;
  assign T324 = T325 | T177;
  assign T325 = T326 | T180;
  assign T326 = T327 | T183;
  assign T327 = T328 | T186;
  assign T328 = T329 | T189;
  assign T329 = T330 | T192;
  assign T330 = T197 | T195;
  assign T331 = T333 & T332;
  assign T332 = R17 < 3'h7;
  assign T333 = T334 ^ 1'h1;
  assign T334 = T335 | T180;
  assign T335 = T336 | T183;
  assign T336 = T337 | T186;
  assign T337 = T338 | T189;
  assign T338 = T339 | T192;
  assign T339 = T197 | T195;

  always @(posedge clk) begin
    if(reset) begin
      R17 <= 3'h0;
    end else if(T19) begin
      R17 <= T0;
    end
  end
endmodule

module RRArbiter_4(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [2:0] io_in_7_bits_payload_master_xact_id,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [2:0] io_in_6_bits_payload_master_xact_id,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [2:0] io_in_5_bits_payload_master_xact_id,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [2:0] io_in_4_bits_payload_master_xact_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [2:0] io_in_3_bits_payload_master_xact_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  reg [2:0] R17;
  wire[2:0] T256;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T38;
  wire T39;
  wire[2:0] T40;
  wire[2:0] T41;
  wire T42;
  wire[2:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire[1:0] T63;
  wire T64;
  wire[1:0] T65;
  wire T66;
  wire T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire T70;
  wire[1:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T30 ? 3'h1 : T2;
  assign T2 = T28 ? 3'h2 : T3;
  assign T3 = T26 ? 3'h3 : T4;
  assign T4 = T24 ? 3'h4 : T5;
  assign T5 = T22 ? 3'h5 : T6;
  assign T6 = T20 ? 3'h6 : T7;
  assign T7 = T15 ? 3'h7 : T8;
  assign T8 = io_in_0_valid ? 3'h0 : T9;
  assign T9 = io_in_1_valid ? 3'h1 : T10;
  assign T10 = io_in_2_valid ? 3'h2 : T11;
  assign T11 = io_in_3_valid ? 3'h3 : T12;
  assign T12 = io_in_4_valid ? 3'h4 : T13;
  assign T13 = io_in_5_valid ? 3'h5 : T14;
  assign T14 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T15 = io_in_7_valid & T16;
  assign T16 = R17 < 3'h7;
  assign T256 = reset ? 3'h0 : T18;
  assign T18 = T19 ? T0 : R17;
  assign T19 = io_out_ready & io_out_valid;
  assign T20 = io_in_6_valid & T21;
  assign T21 = R17 < 3'h6;
  assign T22 = io_in_5_valid & T23;
  assign T23 = R17 < 3'h5;
  assign T24 = io_in_4_valid & T25;
  assign T25 = R17 < 3'h4;
  assign T26 = io_in_3_valid & T27;
  assign T27 = R17 < 3'h3;
  assign T28 = io_in_2_valid & T29;
  assign T29 = R17 < 3'h2;
  assign T30 = io_in_1_valid & T31;
  assign T31 = R17 < 3'h1;
  assign io_out_bits_payload_master_xact_id = T32;
  assign T32 = T46 ? T40 : T33;
  assign T33 = T39 ? T37 : T34;
  assign T34 = T35 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T35 = T36[1'h0:1'h0];
  assign T36 = T0;
  assign T37 = T38 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T38 = T36[1'h0:1'h0];
  assign T39 = T36[1'h1:1'h1];
  assign T40 = T45 ? T43 : T41;
  assign T41 = T42 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T42 = T36[1'h0:1'h0];
  assign T43 = T44 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T44 = T36[1'h0:1'h0];
  assign T45 = T36[1'h1:1'h1];
  assign T46 = T36[2'h2:2'h2];
  assign io_out_bits_header_dst = T47;
  assign T47 = T60 ? T54 : T48;
  assign T48 = T53 ? T51 : T49;
  assign T49 = T50 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T50 = T36[1'h0:1'h0];
  assign T51 = T52 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T52 = T36[1'h0:1'h0];
  assign T53 = T36[1'h1:1'h1];
  assign T54 = T59 ? T57 : T55;
  assign T55 = T56 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T56 = T36[1'h0:1'h0];
  assign T57 = T58 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T58 = T36[1'h0:1'h0];
  assign T59 = T36[1'h1:1'h1];
  assign T60 = T36[2'h2:2'h2];
  assign io_out_bits_header_src = T61;
  assign T61 = T74 ? T68 : T62;
  assign T62 = T67 ? T65 : T63;
  assign T63 = T64 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T64 = T36[1'h0:1'h0];
  assign T65 = T66 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T66 = T36[1'h0:1'h0];
  assign T67 = T36[1'h1:1'h1];
  assign T68 = T73 ? T71 : T69;
  assign T69 = T70 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T70 = T36[1'h0:1'h0];
  assign T71 = T72 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T72 = T36[1'h0:1'h0];
  assign T73 = T36[1'h1:1'h1];
  assign T74 = T36[2'h2:2'h2];
  assign io_out_valid = T75;
  assign T75 = T88 ? T82 : T76;
  assign T76 = T81 ? T79 : T77;
  assign T77 = T78 ? io_in_1_valid : io_in_0_valid;
  assign T78 = T36[1'h0:1'h0];
  assign T79 = T80 ? io_in_3_valid : io_in_2_valid;
  assign T80 = T36[1'h0:1'h0];
  assign T81 = T36[1'h1:1'h1];
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_5_valid : io_in_4_valid;
  assign T84 = T36[1'h0:1'h0];
  assign T85 = T86 ? io_in_7_valid : io_in_6_valid;
  assign T86 = T36[1'h0:1'h0];
  assign T87 = T36[1'h1:1'h1];
  assign T88 = T36[2'h2:2'h2];
  assign io_in_0_ready = T89;
  assign T89 = T90 & io_out_ready;
  assign T90 = T115 | T91;
  assign T91 = T92 ^ 1'h1;
  assign T92 = T95 | T93;
  assign T93 = io_in_7_valid & T94;
  assign T94 = R17 < 3'h7;
  assign T95 = T98 | T96;
  assign T96 = io_in_6_valid & T97;
  assign T97 = R17 < 3'h6;
  assign T98 = T101 | T99;
  assign T99 = io_in_5_valid & T100;
  assign T100 = R17 < 3'h5;
  assign T101 = T104 | T102;
  assign T102 = io_in_4_valid & T103;
  assign T103 = R17 < 3'h4;
  assign T104 = T107 | T105;
  assign T105 = io_in_3_valid & T106;
  assign T106 = R17 < 3'h3;
  assign T107 = T110 | T108;
  assign T108 = io_in_2_valid & T109;
  assign T109 = R17 < 3'h2;
  assign T110 = T113 | T111;
  assign T111 = io_in_1_valid & T112;
  assign T112 = R17 < 3'h1;
  assign T113 = io_in_0_valid & T114;
  assign T114 = R17 < 3'h0;
  assign T115 = R17 < 3'h0;
  assign io_in_1_ready = T116;
  assign T116 = T117 & io_out_ready;
  assign T117 = T127 | T118;
  assign T118 = T119 ^ 1'h1;
  assign T119 = T120 | io_in_0_valid;
  assign T120 = T121 | T93;
  assign T121 = T122 | T96;
  assign T122 = T123 | T99;
  assign T123 = T124 | T102;
  assign T124 = T125 | T105;
  assign T125 = T126 | T108;
  assign T126 = T113 | T111;
  assign T127 = T129 & T128;
  assign T128 = R17 < 3'h1;
  assign T129 = T113 ^ 1'h1;
  assign io_in_2_ready = T130;
  assign T130 = T131 & io_out_ready;
  assign T131 = T142 | T132;
  assign T132 = T133 ^ 1'h1;
  assign T133 = T134 | io_in_1_valid;
  assign T134 = T135 | io_in_0_valid;
  assign T135 = T136 | T93;
  assign T136 = T137 | T96;
  assign T137 = T138 | T99;
  assign T138 = T139 | T102;
  assign T139 = T140 | T105;
  assign T140 = T141 | T108;
  assign T141 = T113 | T111;
  assign T142 = T144 & T143;
  assign T143 = R17 < 3'h2;
  assign T144 = T145 ^ 1'h1;
  assign T145 = T113 | T111;
  assign io_in_3_ready = T146;
  assign T146 = T147 & io_out_ready;
  assign T147 = T159 | T148;
  assign T148 = T149 ^ 1'h1;
  assign T149 = T150 | io_in_2_valid;
  assign T150 = T151 | io_in_1_valid;
  assign T151 = T152 | io_in_0_valid;
  assign T152 = T153 | T93;
  assign T153 = T154 | T96;
  assign T154 = T155 | T99;
  assign T155 = T156 | T102;
  assign T156 = T157 | T105;
  assign T157 = T158 | T108;
  assign T158 = T113 | T111;
  assign T159 = T161 & T160;
  assign T160 = R17 < 3'h3;
  assign T161 = T162 ^ 1'h1;
  assign T162 = T163 | T108;
  assign T163 = T113 | T111;
  assign io_in_4_ready = T164;
  assign T164 = T165 & io_out_ready;
  assign T165 = T178 | T166;
  assign T166 = T167 ^ 1'h1;
  assign T167 = T168 | io_in_3_valid;
  assign T168 = T169 | io_in_2_valid;
  assign T169 = T170 | io_in_1_valid;
  assign T170 = T171 | io_in_0_valid;
  assign T171 = T172 | T93;
  assign T172 = T173 | T96;
  assign T173 = T174 | T99;
  assign T174 = T175 | T102;
  assign T175 = T176 | T105;
  assign T176 = T177 | T108;
  assign T177 = T113 | T111;
  assign T178 = T180 & T179;
  assign T179 = R17 < 3'h4;
  assign T180 = T181 ^ 1'h1;
  assign T181 = T182 | T105;
  assign T182 = T183 | T108;
  assign T183 = T113 | T111;
  assign io_in_5_ready = T184;
  assign T184 = T185 & io_out_ready;
  assign T185 = T199 | T186;
  assign T186 = T187 ^ 1'h1;
  assign T187 = T188 | io_in_4_valid;
  assign T188 = T189 | io_in_3_valid;
  assign T189 = T190 | io_in_2_valid;
  assign T190 = T191 | io_in_1_valid;
  assign T191 = T192 | io_in_0_valid;
  assign T192 = T193 | T93;
  assign T193 = T194 | T96;
  assign T194 = T195 | T99;
  assign T195 = T196 | T102;
  assign T196 = T197 | T105;
  assign T197 = T198 | T108;
  assign T198 = T113 | T111;
  assign T199 = T201 & T200;
  assign T200 = R17 < 3'h5;
  assign T201 = T202 ^ 1'h1;
  assign T202 = T203 | T102;
  assign T203 = T204 | T105;
  assign T204 = T205 | T108;
  assign T205 = T113 | T111;
  assign io_in_6_ready = T206;
  assign T206 = T207 & io_out_ready;
  assign T207 = T222 | T208;
  assign T208 = T209 ^ 1'h1;
  assign T209 = T210 | io_in_5_valid;
  assign T210 = T211 | io_in_4_valid;
  assign T211 = T212 | io_in_3_valid;
  assign T212 = T213 | io_in_2_valid;
  assign T213 = T214 | io_in_1_valid;
  assign T214 = T215 | io_in_0_valid;
  assign T215 = T216 | T93;
  assign T216 = T217 | T96;
  assign T217 = T218 | T99;
  assign T218 = T219 | T102;
  assign T219 = T220 | T105;
  assign T220 = T221 | T108;
  assign T221 = T113 | T111;
  assign T222 = T224 & T223;
  assign T223 = R17 < 3'h6;
  assign T224 = T225 ^ 1'h1;
  assign T225 = T226 | T99;
  assign T226 = T227 | T102;
  assign T227 = T228 | T105;
  assign T228 = T229 | T108;
  assign T229 = T113 | T111;
  assign io_in_7_ready = T230;
  assign T230 = T231 & io_out_ready;
  assign T231 = T247 | T232;
  assign T232 = T233 ^ 1'h1;
  assign T233 = T234 | io_in_6_valid;
  assign T234 = T235 | io_in_5_valid;
  assign T235 = T236 | io_in_4_valid;
  assign T236 = T237 | io_in_3_valid;
  assign T237 = T238 | io_in_2_valid;
  assign T238 = T239 | io_in_1_valid;
  assign T239 = T240 | io_in_0_valid;
  assign T240 = T241 | T93;
  assign T241 = T242 | T96;
  assign T242 = T243 | T99;
  assign T243 = T244 | T102;
  assign T244 = T245 | T105;
  assign T245 = T246 | T108;
  assign T246 = T113 | T111;
  assign T247 = T249 & T248;
  assign T248 = R17 < 3'h7;
  assign T249 = T250 ^ 1'h1;
  assign T250 = T251 | T96;
  assign T251 = T252 | T99;
  assign T252 = T253 | T102;
  assign T253 = T254 | T105;
  assign T254 = T255 | T108;
  assign T255 = T113 | T111;

  always @(posedge clk) begin
    if(reset) begin
      R17 <= 3'h0;
    end else if(T19) begin
      R17 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatPassesId(input clk, input reset,
    output io_in_7_acquire_ready,
    input  io_in_7_acquire_valid,
    input [1:0] io_in_7_acquire_bits_header_src,
    input [1:0] io_in_7_acquire_bits_header_dst,
    input [25:0] io_in_7_acquire_bits_payload_addr,
    input [1:0] io_in_7_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_7_acquire_bits_payload_data,
    input [2:0] io_in_7_acquire_bits_payload_a_type,
    input [5:0] io_in_7_acquire_bits_payload_write_mask,
    input [2:0] io_in_7_acquire_bits_payload_subword_addr,
    input [3:0] io_in_7_acquire_bits_payload_atomic_opcode,
    input  io_in_7_grant_ready,
    output io_in_7_grant_valid,
    output[1:0] io_in_7_grant_bits_header_src,
    output[1:0] io_in_7_grant_bits_header_dst,
    output[511:0] io_in_7_grant_bits_payload_data,
    output[1:0] io_in_7_grant_bits_payload_client_xact_id,
    output[2:0] io_in_7_grant_bits_payload_master_xact_id,
    output[3:0] io_in_7_grant_bits_payload_g_type,
    output io_in_7_finish_ready,
    input  io_in_7_finish_valid,
    input [1:0] io_in_7_finish_bits_header_src,
    input [1:0] io_in_7_finish_bits_header_dst,
    input [2:0] io_in_7_finish_bits_payload_master_xact_id,
    output io_in_6_acquire_ready,
    input  io_in_6_acquire_valid,
    input [1:0] io_in_6_acquire_bits_header_src,
    input [1:0] io_in_6_acquire_bits_header_dst,
    input [25:0] io_in_6_acquire_bits_payload_addr,
    input [1:0] io_in_6_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_6_acquire_bits_payload_data,
    input [2:0] io_in_6_acquire_bits_payload_a_type,
    input [5:0] io_in_6_acquire_bits_payload_write_mask,
    input [2:0] io_in_6_acquire_bits_payload_subword_addr,
    input [3:0] io_in_6_acquire_bits_payload_atomic_opcode,
    input  io_in_6_grant_ready,
    output io_in_6_grant_valid,
    output[1:0] io_in_6_grant_bits_header_src,
    output[1:0] io_in_6_grant_bits_header_dst,
    output[511:0] io_in_6_grant_bits_payload_data,
    output[1:0] io_in_6_grant_bits_payload_client_xact_id,
    output[2:0] io_in_6_grant_bits_payload_master_xact_id,
    output[3:0] io_in_6_grant_bits_payload_g_type,
    output io_in_6_finish_ready,
    input  io_in_6_finish_valid,
    input [1:0] io_in_6_finish_bits_header_src,
    input [1:0] io_in_6_finish_bits_header_dst,
    input [2:0] io_in_6_finish_bits_payload_master_xact_id,
    output io_in_5_acquire_ready,
    input  io_in_5_acquire_valid,
    input [1:0] io_in_5_acquire_bits_header_src,
    input [1:0] io_in_5_acquire_bits_header_dst,
    input [25:0] io_in_5_acquire_bits_payload_addr,
    input [1:0] io_in_5_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_5_acquire_bits_payload_data,
    input [2:0] io_in_5_acquire_bits_payload_a_type,
    input [5:0] io_in_5_acquire_bits_payload_write_mask,
    input [2:0] io_in_5_acquire_bits_payload_subword_addr,
    input [3:0] io_in_5_acquire_bits_payload_atomic_opcode,
    input  io_in_5_grant_ready,
    output io_in_5_grant_valid,
    output[1:0] io_in_5_grant_bits_header_src,
    output[1:0] io_in_5_grant_bits_header_dst,
    output[511:0] io_in_5_grant_bits_payload_data,
    output[1:0] io_in_5_grant_bits_payload_client_xact_id,
    output[2:0] io_in_5_grant_bits_payload_master_xact_id,
    output[3:0] io_in_5_grant_bits_payload_g_type,
    output io_in_5_finish_ready,
    input  io_in_5_finish_valid,
    input [1:0] io_in_5_finish_bits_header_src,
    input [1:0] io_in_5_finish_bits_header_dst,
    input [2:0] io_in_5_finish_bits_payload_master_xact_id,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [1:0] io_in_4_acquire_bits_header_src,
    input [1:0] io_in_4_acquire_bits_header_dst,
    input [25:0] io_in_4_acquire_bits_payload_addr,
    input [1:0] io_in_4_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_4_acquire_bits_payload_data,
    input [2:0] io_in_4_acquire_bits_payload_a_type,
    input [5:0] io_in_4_acquire_bits_payload_write_mask,
    input [2:0] io_in_4_acquire_bits_payload_subword_addr,
    input [3:0] io_in_4_acquire_bits_payload_atomic_opcode,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_header_src,
    output[1:0] io_in_4_grant_bits_header_dst,
    output[511:0] io_in_4_grant_bits_payload_data,
    output[1:0] io_in_4_grant_bits_payload_client_xact_id,
    output[2:0] io_in_4_grant_bits_payload_master_xact_id,
    output[3:0] io_in_4_grant_bits_payload_g_type,
    output io_in_4_finish_ready,
    input  io_in_4_finish_valid,
    input [1:0] io_in_4_finish_bits_header_src,
    input [1:0] io_in_4_finish_bits_header_dst,
    input [2:0] io_in_4_finish_bits_payload_master_xact_id,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [1:0] io_in_3_acquire_bits_header_src,
    input [1:0] io_in_3_acquire_bits_header_dst,
    input [25:0] io_in_3_acquire_bits_payload_addr,
    input [1:0] io_in_3_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_3_acquire_bits_payload_data,
    input [2:0] io_in_3_acquire_bits_payload_a_type,
    input [5:0] io_in_3_acquire_bits_payload_write_mask,
    input [2:0] io_in_3_acquire_bits_payload_subword_addr,
    input [3:0] io_in_3_acquire_bits_payload_atomic_opcode,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_header_src,
    output[1:0] io_in_3_grant_bits_header_dst,
    output[511:0] io_in_3_grant_bits_payload_data,
    output[1:0] io_in_3_grant_bits_payload_client_xact_id,
    output[2:0] io_in_3_grant_bits_payload_master_xact_id,
    output[3:0] io_in_3_grant_bits_payload_g_type,
    output io_in_3_finish_ready,
    input  io_in_3_finish_valid,
    input [1:0] io_in_3_finish_bits_header_src,
    input [1:0] io_in_3_finish_bits_header_dst,
    input [2:0] io_in_3_finish_bits_payload_master_xact_id,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [1:0] io_in_2_acquire_bits_header_src,
    input [1:0] io_in_2_acquire_bits_header_dst,
    input [25:0] io_in_2_acquire_bits_payload_addr,
    input [1:0] io_in_2_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_2_acquire_bits_payload_data,
    input [2:0] io_in_2_acquire_bits_payload_a_type,
    input [5:0] io_in_2_acquire_bits_payload_write_mask,
    input [2:0] io_in_2_acquire_bits_payload_subword_addr,
    input [3:0] io_in_2_acquire_bits_payload_atomic_opcode,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_header_src,
    output[1:0] io_in_2_grant_bits_header_dst,
    output[511:0] io_in_2_grant_bits_payload_data,
    output[1:0] io_in_2_grant_bits_payload_client_xact_id,
    output[2:0] io_in_2_grant_bits_payload_master_xact_id,
    output[3:0] io_in_2_grant_bits_payload_g_type,
    output io_in_2_finish_ready,
    input  io_in_2_finish_valid,
    input [1:0] io_in_2_finish_bits_header_src,
    input [1:0] io_in_2_finish_bits_header_dst,
    input [2:0] io_in_2_finish_bits_payload_master_xact_id,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [1:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_1_acquire_bits_payload_data,
    input [2:0] io_in_1_acquire_bits_payload_a_type,
    input [5:0] io_in_1_acquire_bits_payload_write_mask,
    input [2:0] io_in_1_acquire_bits_payload_subword_addr,
    input [3:0] io_in_1_acquire_bits_payload_atomic_opcode,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[511:0] io_in_1_grant_bits_payload_data,
    output[1:0] io_in_1_grant_bits_payload_client_xact_id,
    output[2:0] io_in_1_grant_bits_payload_master_xact_id,
    output[3:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input [2:0] io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [1:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_0_acquire_bits_payload_data,
    input [2:0] io_in_0_acquire_bits_payload_a_type,
    input [5:0] io_in_0_acquire_bits_payload_write_mask,
    input [2:0] io_in_0_acquire_bits_payload_subword_addr,
    input [3:0] io_in_0_acquire_bits_payload_atomic_opcode,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[511:0] io_in_0_grant_bits_payload_data,
    output[1:0] io_in_0_grant_bits_payload_client_xact_id,
    output[2:0] io_in_0_grant_bits_payload_master_xact_id,
    output[3:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input [2:0] io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[1:0] io_out_acquire_bits_payload_client_xact_id,
    output[511:0] io_out_acquire_bits_payload_data,
    output[2:0] io_out_acquire_bits_payload_a_type,
    output[5:0] io_out_acquire_bits_payload_write_mask,
    output[2:0] io_out_acquire_bits_payload_subword_addr,
    output[3:0] io_out_acquire_bits_payload_atomic_opcode,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [511:0] io_out_grant_bits_payload_data,
    input [1:0] io_out_grant_bits_payload_client_xact_id,
    input [2:0] io_out_grant_bits_payload_master_xact_id,
    input [3:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[2:0] io_out_finish_bits_payload_master_xact_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] T24;
  wire T13;
  wire[2:0] T25;
  wire T14;
  wire[2:0] T26;
  wire T15;
  wire[2:0] T27;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire RRArbiter_2_io_in_7_ready;
  wire RRArbiter_2_io_in_6_ready;
  wire RRArbiter_2_io_in_5_ready;
  wire RRArbiter_2_io_in_4_ready;
  wire RRArbiter_2_io_in_3_ready;
  wire RRArbiter_2_io_in_2_ready;
  wire RRArbiter_2_io_in_1_ready;
  wire RRArbiter_2_io_in_0_ready;
  wire RRArbiter_2_io_out_valid;
  wire[1:0] RRArbiter_2_io_out_bits_header_src;
  wire[1:0] RRArbiter_2_io_out_bits_header_dst;
  wire[25:0] RRArbiter_2_io_out_bits_payload_addr;
  wire[1:0] RRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[511:0] RRArbiter_2_io_out_bits_payload_data;
  wire[2:0] RRArbiter_2_io_out_bits_payload_a_type;
  wire[5:0] RRArbiter_2_io_out_bits_payload_write_mask;
  wire[2:0] RRArbiter_2_io_out_bits_payload_subword_addr;
  wire[3:0] RRArbiter_2_io_out_bits_payload_atomic_opcode;
  wire RRArbiter_3_io_in_7_ready;
  wire RRArbiter_3_io_in_6_ready;
  wire RRArbiter_3_io_in_5_ready;
  wire RRArbiter_3_io_in_4_ready;
  wire RRArbiter_3_io_in_3_ready;
  wire RRArbiter_3_io_in_2_ready;
  wire RRArbiter_3_io_in_1_ready;
  wire RRArbiter_3_io_in_0_ready;
  wire RRArbiter_3_io_out_valid;
  wire[1:0] RRArbiter_3_io_out_bits_header_src;
  wire[1:0] RRArbiter_3_io_out_bits_header_dst;
  wire[2:0] RRArbiter_3_io_out_bits_payload_master_xact_id;


  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_3_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_3_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_3_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_3_io_out_valid;
  assign io_out_grant_ready = T0;
  assign T0 = T15 ? io_in_7_grant_ready : T1;
  assign T1 = T14 ? io_in_6_grant_ready : T2;
  assign T2 = T13 ? io_in_5_grant_ready : T3;
  assign T3 = T12 ? io_in_4_grant_ready : T4;
  assign T4 = T11 ? io_in_3_grant_ready : T5;
  assign T5 = T10 ? io_in_2_grant_ready : T6;
  assign T6 = T9 ? io_in_1_grant_ready : T7;
  assign T7 = T8 ? io_in_0_grant_ready : 1'h0;
  assign T8 = io_out_grant_bits_payload_client_xact_id == 2'h0;
  assign T9 = io_out_grant_bits_payload_client_xact_id == 2'h1;
  assign T10 = io_out_grant_bits_payload_client_xact_id == 2'h2;
  assign T11 = io_out_grant_bits_payload_client_xact_id == 2'h3;
  assign T12 = T24 == 3'h4;
  assign T24 = {1'h0, io_out_grant_bits_payload_client_xact_id};
  assign T13 = T25 == 3'h5;
  assign T25 = {1'h0, io_out_grant_bits_payload_client_xact_id};
  assign T14 = T26 == 3'h6;
  assign T26 = {1'h0, io_out_grant_bits_payload_client_xact_id};
  assign T15 = T27 == 3'h7;
  assign T27 = {1'h0, io_out_grant_bits_payload_client_xact_id};
  assign io_out_acquire_bits_payload_atomic_opcode = RRArbiter_2_io_out_bits_payload_atomic_opcode;
  assign io_out_acquire_bits_payload_subword_addr = RRArbiter_2_io_out_bits_payload_subword_addr;
  assign io_out_acquire_bits_payload_write_mask = RRArbiter_2_io_out_bits_payload_write_mask;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_2_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_data = RRArbiter_2_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_2_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_2_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_2_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_2_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_3_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T16;
  assign T16 = T8 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_2_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_3_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T17;
  assign T17 = T9 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_2_io_in_1_ready;
  assign io_in_2_finish_ready = RRArbiter_3_io_in_2_ready;
  assign io_in_2_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_2_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_2_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_2_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_2_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_2_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_2_grant_valid = T18;
  assign T18 = T10 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = RRArbiter_2_io_in_2_ready;
  assign io_in_3_finish_ready = RRArbiter_3_io_in_3_ready;
  assign io_in_3_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_3_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_3_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_3_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_3_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_3_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_3_grant_valid = T19;
  assign T19 = T11 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = RRArbiter_2_io_in_3_ready;
  assign io_in_4_finish_ready = RRArbiter_3_io_in_4_ready;
  assign io_in_4_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_4_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_4_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_4_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_4_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_4_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_4_grant_valid = T20;
  assign T20 = T12 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = RRArbiter_2_io_in_4_ready;
  assign io_in_5_finish_ready = RRArbiter_3_io_in_5_ready;
  assign io_in_5_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_5_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_5_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_5_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_5_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_5_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_5_grant_valid = T21;
  assign T21 = T13 ? io_out_grant_valid : 1'h0;
  assign io_in_5_acquire_ready = RRArbiter_2_io_in_5_ready;
  assign io_in_6_finish_ready = RRArbiter_3_io_in_6_ready;
  assign io_in_6_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_6_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_6_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_6_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_6_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_6_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_6_grant_valid = T22;
  assign T22 = T14 ? io_out_grant_valid : 1'h0;
  assign io_in_6_acquire_ready = RRArbiter_2_io_in_6_ready;
  assign io_in_7_finish_ready = RRArbiter_3_io_in_7_ready;
  assign io_in_7_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_7_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_7_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_7_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_7_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_7_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_7_grant_valid = T23;
  assign T23 = T15 ? io_out_grant_valid : 1'h0;
  assign io_in_7_acquire_ready = RRArbiter_2_io_in_7_ready;
  RRArbiter_3 RRArbiter_2(.clk(clk), .reset(reset),
       .io_in_7_ready( RRArbiter_2_io_in_7_ready ),
       .io_in_7_valid( io_in_7_acquire_valid ),
       .io_in_7_bits_header_src( io_in_7_acquire_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_acquire_bits_header_dst ),
       .io_in_7_bits_payload_addr( io_in_7_acquire_bits_payload_addr ),
       .io_in_7_bits_payload_client_xact_id( io_in_7_acquire_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_data( io_in_7_acquire_bits_payload_data ),
       .io_in_7_bits_payload_a_type( io_in_7_acquire_bits_payload_a_type ),
       .io_in_7_bits_payload_write_mask( io_in_7_acquire_bits_payload_write_mask ),
       .io_in_7_bits_payload_subword_addr( io_in_7_acquire_bits_payload_subword_addr ),
       .io_in_7_bits_payload_atomic_opcode( io_in_7_acquire_bits_payload_atomic_opcode ),
       .io_in_6_ready( RRArbiter_2_io_in_6_ready ),
       .io_in_6_valid( io_in_6_acquire_valid ),
       .io_in_6_bits_header_src( io_in_6_acquire_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_acquire_bits_header_dst ),
       .io_in_6_bits_payload_addr( io_in_6_acquire_bits_payload_addr ),
       .io_in_6_bits_payload_client_xact_id( io_in_6_acquire_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_data( io_in_6_acquire_bits_payload_data ),
       .io_in_6_bits_payload_a_type( io_in_6_acquire_bits_payload_a_type ),
       .io_in_6_bits_payload_write_mask( io_in_6_acquire_bits_payload_write_mask ),
       .io_in_6_bits_payload_subword_addr( io_in_6_acquire_bits_payload_subword_addr ),
       .io_in_6_bits_payload_atomic_opcode( io_in_6_acquire_bits_payload_atomic_opcode ),
       .io_in_5_ready( RRArbiter_2_io_in_5_ready ),
       .io_in_5_valid( io_in_5_acquire_valid ),
       .io_in_5_bits_header_src( io_in_5_acquire_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_acquire_bits_header_dst ),
       .io_in_5_bits_payload_addr( io_in_5_acquire_bits_payload_addr ),
       .io_in_5_bits_payload_client_xact_id( io_in_5_acquire_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_data( io_in_5_acquire_bits_payload_data ),
       .io_in_5_bits_payload_a_type( io_in_5_acquire_bits_payload_a_type ),
       .io_in_5_bits_payload_write_mask( io_in_5_acquire_bits_payload_write_mask ),
       .io_in_5_bits_payload_subword_addr( io_in_5_acquire_bits_payload_subword_addr ),
       .io_in_5_bits_payload_atomic_opcode( io_in_5_acquire_bits_payload_atomic_opcode ),
       .io_in_4_ready( RRArbiter_2_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_header_src( io_in_4_acquire_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_acquire_bits_header_dst ),
       .io_in_4_bits_payload_addr( io_in_4_acquire_bits_payload_addr ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_acquire_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_data( io_in_4_acquire_bits_payload_data ),
       .io_in_4_bits_payload_a_type( io_in_4_acquire_bits_payload_a_type ),
       .io_in_4_bits_payload_write_mask( io_in_4_acquire_bits_payload_write_mask ),
       .io_in_4_bits_payload_subword_addr( io_in_4_acquire_bits_payload_subword_addr ),
       .io_in_4_bits_payload_atomic_opcode( io_in_4_acquire_bits_payload_atomic_opcode ),
       .io_in_3_ready( RRArbiter_2_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_header_src( io_in_3_acquire_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_acquire_bits_header_dst ),
       .io_in_3_bits_payload_addr( io_in_3_acquire_bits_payload_addr ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_acquire_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_data( io_in_3_acquire_bits_payload_data ),
       .io_in_3_bits_payload_a_type( io_in_3_acquire_bits_payload_a_type ),
       .io_in_3_bits_payload_write_mask( io_in_3_acquire_bits_payload_write_mask ),
       .io_in_3_bits_payload_subword_addr( io_in_3_acquire_bits_payload_subword_addr ),
       .io_in_3_bits_payload_atomic_opcode( io_in_3_acquire_bits_payload_atomic_opcode ),
       .io_in_2_ready( RRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_header_src( io_in_2_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_acquire_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_acquire_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_acquire_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_acquire_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_acquire_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_acquire_bits_payload_atomic_opcode ),
       .io_in_1_ready( RRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_acquire_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_acquire_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_acquire_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_acquire_bits_payload_atomic_opcode ),
       .io_in_0_ready( RRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_acquire_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_acquire_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_acquire_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_acquire_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( RRArbiter_2_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( RRArbiter_2_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( RRArbiter_2_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( RRArbiter_2_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  RRArbiter_4 RRArbiter_3(.clk(clk), .reset(reset),
       .io_in_7_ready( RRArbiter_3_io_in_7_ready ),
       .io_in_7_valid( io_in_7_finish_valid ),
       .io_in_7_bits_header_src( io_in_7_finish_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_finish_bits_header_dst ),
       .io_in_7_bits_payload_master_xact_id( io_in_7_finish_bits_payload_master_xact_id ),
       .io_in_6_ready( RRArbiter_3_io_in_6_ready ),
       .io_in_6_valid( io_in_6_finish_valid ),
       .io_in_6_bits_header_src( io_in_6_finish_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_finish_bits_header_dst ),
       .io_in_6_bits_payload_master_xact_id( io_in_6_finish_bits_payload_master_xact_id ),
       .io_in_5_ready( RRArbiter_3_io_in_5_ready ),
       .io_in_5_valid( io_in_5_finish_valid ),
       .io_in_5_bits_header_src( io_in_5_finish_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_finish_bits_header_dst ),
       .io_in_5_bits_payload_master_xact_id( io_in_5_finish_bits_payload_master_xact_id ),
       .io_in_4_ready( RRArbiter_3_io_in_4_ready ),
       .io_in_4_valid( io_in_4_finish_valid ),
       .io_in_4_bits_header_src( io_in_4_finish_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_finish_bits_header_dst ),
       .io_in_4_bits_payload_master_xact_id( io_in_4_finish_bits_payload_master_xact_id ),
       .io_in_3_ready( RRArbiter_3_io_in_3_ready ),
       .io_in_3_valid( io_in_3_finish_valid ),
       .io_in_3_bits_header_src( io_in_3_finish_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_finish_bits_header_dst ),
       .io_in_3_bits_payload_master_xact_id( io_in_3_finish_bits_payload_master_xact_id ),
       .io_in_2_ready( RRArbiter_3_io_in_2_ready ),
       .io_in_2_valid( io_in_2_finish_valid ),
       .io_in_2_bits_header_src( io_in_2_finish_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_finish_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_finish_bits_payload_master_xact_id ),
       .io_in_1_ready( RRArbiter_3_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_3_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_3_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_3_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_3_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_3_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module L2CoherenceAgent(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    output[1:0] io_outer_acquire_bits_header_dst,
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    output io_outer_finish_valid,
    output[1:0] io_outer_finish_bits_header_src,
    output[1:0] io_outer_finish_bits_header_dst,
    output[2:0] io_outer_finish_bits_payload_master_xact_id,
    input  io_incoherent_1,
    input  io_incoherent_0
);

  wire T30;
  wire T31;
  wire any_acquire_conflict;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire[2:0] release_idx;
  wire voluntary;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire T40;
  wire T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire T55;
  wire T56;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire VoluntaryReleaseTracker_io_inner_acquire_ready;
  wire VoluntaryReleaseTracker_io_inner_grant_valid;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_src;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_dst;
  wire[511:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_data;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type;
  wire VoluntaryReleaseTracker_io_inner_probe_valid;
  wire VoluntaryReleaseTracker_io_inner_release_ready;
  wire VoluntaryReleaseTracker_io_outer_acquire_valid;
  wire[1:0] VoluntaryReleaseTracker_io_outer_acquire_bits_header_src;
  wire[25:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr;
  wire[1:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type;
  wire[5:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode;
  wire VoluntaryReleaseTracker_io_outer_grant_ready;
  wire VoluntaryReleaseTracker_io_has_acquire_conflict;
  wire AcquireTracker_0_io_inner_acquire_ready;
  wire AcquireTracker_0_io_inner_grant_valid;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_0_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_0_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_0_io_inner_probe_valid;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_0_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_0_io_inner_release_ready;
  wire AcquireTracker_0_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_0_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_0_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_0_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_0_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_0_io_outer_grant_ready;
  wire AcquireTracker_0_io_has_acquire_conflict;
  wire AcquireTracker_1_io_inner_acquire_ready;
  wire AcquireTracker_1_io_inner_grant_valid;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_1_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_1_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_1_io_inner_probe_valid;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_1_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_1_io_inner_release_ready;
  wire AcquireTracker_1_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_1_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_1_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_1_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_1_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_1_io_outer_grant_ready;
  wire AcquireTracker_1_io_has_acquire_conflict;
  wire AcquireTracker_2_io_inner_acquire_ready;
  wire AcquireTracker_2_io_inner_grant_valid;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_2_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_2_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_2_io_inner_probe_valid;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_2_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_2_io_inner_release_ready;
  wire AcquireTracker_2_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_2_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_2_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_2_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_2_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_2_io_outer_grant_ready;
  wire AcquireTracker_2_io_has_acquire_conflict;
  wire AcquireTracker_3_io_inner_acquire_ready;
  wire AcquireTracker_3_io_inner_grant_valid;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_3_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_3_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_3_io_inner_probe_valid;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_3_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_3_io_inner_release_ready;
  wire AcquireTracker_3_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_3_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_3_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_3_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_3_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_3_io_outer_grant_ready;
  wire AcquireTracker_3_io_has_acquire_conflict;
  wire AcquireTracker_4_io_inner_acquire_ready;
  wire AcquireTracker_4_io_inner_grant_valid;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_4_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_4_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_4_io_inner_probe_valid;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_4_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_4_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_4_io_inner_release_ready;
  wire AcquireTracker_4_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_4_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_4_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_4_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_4_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_4_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_4_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_4_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_4_io_outer_grant_ready;
  wire AcquireTracker_4_io_has_acquire_conflict;
  wire AcquireTracker_5_io_inner_acquire_ready;
  wire AcquireTracker_5_io_inner_grant_valid;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_5_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_5_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_5_io_inner_probe_valid;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_5_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_5_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_5_io_inner_release_ready;
  wire AcquireTracker_5_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_5_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_5_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_5_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_5_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_5_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_5_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_5_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_5_io_outer_grant_ready;
  wire AcquireTracker_5_io_has_acquire_conflict;
  wire AcquireTracker_6_io_inner_acquire_ready;
  wire AcquireTracker_6_io_inner_grant_valid;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_src;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_dst;
  wire[511:0] AcquireTracker_6_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] AcquireTracker_6_io_inner_grant_bits_payload_g_type;
  wire AcquireTracker_6_io_inner_probe_valid;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_src;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_dst;
  wire[25:0] AcquireTracker_6_io_inner_probe_bits_payload_addr;
  wire[2:0] AcquireTracker_6_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_payload_p_type;
  wire AcquireTracker_6_io_inner_release_ready;
  wire AcquireTracker_6_io_outer_acquire_valid;
  wire[1:0] AcquireTracker_6_io_outer_acquire_bits_header_src;
  wire[25:0] AcquireTracker_6_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_6_io_outer_acquire_bits_payload_data;
  wire[2:0] AcquireTracker_6_io_outer_acquire_bits_payload_a_type;
  wire[5:0] AcquireTracker_6_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_6_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] AcquireTracker_6_io_outer_acquire_bits_payload_atomic_opcode;
  wire AcquireTracker_6_io_outer_grant_ready;
  wire AcquireTracker_6_io_has_acquire_conflict;
  wire alloc_arb_io_in_7_ready;
  wire alloc_arb_io_in_6_ready;
  wire alloc_arb_io_in_5_ready;
  wire alloc_arb_io_in_4_ready;
  wire alloc_arb_io_in_3_ready;
  wire alloc_arb_io_in_2_ready;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire probe_arb_io_in_7_ready;
  wire probe_arb_io_in_6_ready;
  wire probe_arb_io_in_5_ready;
  wire probe_arb_io_in_4_ready;
  wire probe_arb_io_in_3_ready;
  wire probe_arb_io_in_2_ready;
  wire probe_arb_io_in_1_ready;
  wire probe_arb_io_in_0_ready;
  wire probe_arb_io_out_valid;
  wire[1:0] probe_arb_io_out_bits_header_src;
  wire[1:0] probe_arb_io_out_bits_header_dst;
  wire[25:0] probe_arb_io_out_bits_payload_addr;
  wire[2:0] probe_arb_io_out_bits_payload_master_xact_id;
  wire[1:0] probe_arb_io_out_bits_payload_p_type;
  wire grant_arb_io_in_7_ready;
  wire grant_arb_io_in_6_ready;
  wire grant_arb_io_in_5_ready;
  wire grant_arb_io_in_4_ready;
  wire grant_arb_io_in_3_ready;
  wire grant_arb_io_in_2_ready;
  wire grant_arb_io_in_1_ready;
  wire grant_arb_io_in_0_ready;
  wire grant_arb_io_out_valid;
  wire[1:0] grant_arb_io_out_bits_header_src;
  wire[1:0] grant_arb_io_out_bits_header_dst;
  wire[511:0] grant_arb_io_out_bits_payload_data;
  wire[1:0] grant_arb_io_out_bits_payload_client_xact_id;
  wire[2:0] grant_arb_io_out_bits_payload_master_xact_id;
  wire[3:0] grant_arb_io_out_bits_payload_g_type;
  wire outer_arb_io_in_7_acquire_ready;
  wire outer_arb_io_in_7_grant_valid;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_7_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_7_grant_bits_payload_client_xact_id;
  wire[2:0] outer_arb_io_in_7_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_7_grant_bits_payload_g_type;
  wire outer_arb_io_in_7_finish_ready;
  wire outer_arb_io_in_6_acquire_ready;
  wire outer_arb_io_in_6_grant_valid;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_6_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_6_grant_bits_payload_client_xact_id;
  wire[2:0] outer_arb_io_in_6_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_6_grant_bits_payload_g_type;
  wire outer_arb_io_in_6_finish_ready;
  wire outer_arb_io_in_5_acquire_ready;
  wire outer_arb_io_in_5_grant_valid;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_5_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_5_grant_bits_payload_client_xact_id;
  wire[2:0] outer_arb_io_in_5_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_5_grant_bits_payload_g_type;
  wire outer_arb_io_in_5_finish_ready;
  wire outer_arb_io_in_4_acquire_ready;
  wire outer_arb_io_in_4_grant_valid;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_4_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_4_grant_bits_payload_client_xact_id;
  wire[2:0] outer_arb_io_in_4_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_4_grant_bits_payload_g_type;
  wire outer_arb_io_in_4_finish_ready;
  wire outer_arb_io_in_3_acquire_ready;
  wire outer_arb_io_in_3_grant_valid;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_3_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_3_grant_bits_payload_client_xact_id;
  wire[2:0] outer_arb_io_in_3_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_3_grant_bits_payload_g_type;
  wire outer_arb_io_in_3_finish_ready;
  wire outer_arb_io_in_2_acquire_ready;
  wire outer_arb_io_in_2_grant_valid;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_2_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_2_grant_bits_payload_client_xact_id;
  wire[2:0] outer_arb_io_in_2_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_2_grant_bits_payload_g_type;
  wire outer_arb_io_in_2_finish_ready;
  wire outer_arb_io_in_1_acquire_ready;
  wire outer_arb_io_in_1_grant_valid;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_1_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_1_grant_bits_payload_client_xact_id;
  wire[2:0] outer_arb_io_in_1_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_1_grant_bits_payload_g_type;
  wire outer_arb_io_in_1_finish_ready;
  wire outer_arb_io_in_0_acquire_ready;
  wire outer_arb_io_in_0_grant_valid;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_src;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_dst;
  wire[511:0] outer_arb_io_in_0_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_0_grant_bits_payload_client_xact_id;
  wire[2:0] outer_arb_io_in_0_grant_bits_payload_master_xact_id;
  wire[3:0] outer_arb_io_in_0_grant_bits_payload_g_type;
  wire outer_arb_io_in_0_finish_ready;
  wire outer_arb_io_out_acquire_valid;
  wire[1:0] outer_arb_io_out_acquire_bits_header_src;
  wire[1:0] outer_arb_io_out_acquire_bits_header_dst;
  wire[25:0] outer_arb_io_out_acquire_bits_payload_addr;
  wire[1:0] outer_arb_io_out_acquire_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_out_acquire_bits_payload_data;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_a_type;
  wire[5:0] outer_arb_io_out_acquire_bits_payload_write_mask;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_subword_addr;
  wire[3:0] outer_arb_io_out_acquire_bits_payload_atomic_opcode;
  wire outer_arb_io_out_grant_ready;
  wire outer_arb_io_out_finish_valid;
  wire[1:0] outer_arb_io_out_finish_bits_header_src;
  wire[1:0] outer_arb_io_out_finish_bits_header_dst;
  wire[2:0] outer_arb_io_out_finish_bits_payload_master_xact_id;


  assign T30 = io_inner_acquire_valid & T31;
  assign T31 = any_acquire_conflict ^ 1'h1;
  assign any_acquire_conflict = T17 | AcquireTracker_6_io_has_acquire_conflict;
  assign T17 = T18 | AcquireTracker_5_io_has_acquire_conflict;
  assign T18 = T19 | AcquireTracker_4_io_has_acquire_conflict;
  assign T19 = T20 | AcquireTracker_3_io_has_acquire_conflict;
  assign T20 = T21 | AcquireTracker_2_io_has_acquire_conflict;
  assign T21 = T22 | AcquireTracker_1_io_has_acquire_conflict;
  assign T22 = VoluntaryReleaseTracker_io_has_acquire_conflict | AcquireTracker_0_io_has_acquire_conflict;
  assign T32 = T33;
  assign T33 = {io_incoherent_1, io_incoherent_0};
  assign T34 = io_inner_release_valid & T35;
  assign T35 = release_idx == 3'h7;
  assign release_idx = voluntary ? 3'h0 : io_inner_release_bits_payload_master_xact_id;
  assign voluntary = io_inner_release_bits_payload_r_type == 3'h0;
  assign T36 = T33;
  assign T37 = io_inner_release_valid & T38;
  assign T38 = release_idx == 3'h6;
  assign T39 = T33;
  assign T40 = io_inner_release_valid & T41;
  assign T41 = release_idx == 3'h5;
  assign T42 = T33;
  assign T43 = io_inner_release_valid & T44;
  assign T44 = release_idx == 3'h4;
  assign T45 = T33;
  assign T46 = io_inner_release_valid & T47;
  assign T47 = release_idx == 3'h3;
  assign T48 = T33;
  assign T49 = io_inner_release_valid & T50;
  assign T50 = release_idx == 3'h2;
  assign T51 = T33;
  assign T52 = io_inner_release_valid & T53;
  assign T53 = release_idx == 3'h1;
  assign T54 = T33;
  assign T55 = io_inner_release_valid & T56;
  assign T56 = release_idx == 3'h0;
  assign io_outer_finish_bits_payload_master_xact_id = outer_arb_io_out_finish_bits_payload_master_xact_id;
  assign io_outer_finish_bits_header_dst = outer_arb_io_out_finish_bits_header_dst;
  assign io_outer_finish_bits_header_src = outer_arb_io_out_finish_bits_header_src;
  assign io_outer_finish_valid = outer_arb_io_out_finish_valid;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = outer_arb_io_out_acquire_bits_payload_atomic_opcode;
  assign io_outer_acquire_bits_payload_subword_addr = outer_arb_io_out_acquire_bits_payload_subword_addr;
  assign io_outer_acquire_bits_payload_write_mask = outer_arb_io_out_acquire_bits_payload_write_mask;
  assign io_outer_acquire_bits_payload_a_type = outer_arb_io_out_acquire_bits_payload_a_type;
  assign io_outer_acquire_bits_payload_data = outer_arb_io_out_acquire_bits_payload_data;
  assign io_outer_acquire_bits_payload_client_xact_id = outer_arb_io_out_acquire_bits_payload_client_xact_id;
  assign io_outer_acquire_bits_payload_addr = outer_arb_io_out_acquire_bits_payload_addr;
  assign io_outer_acquire_bits_header_dst = outer_arb_io_out_acquire_bits_header_dst;
  assign io_outer_acquire_bits_header_src = outer_arb_io_out_acquire_bits_header_src;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T0;
  assign T0 = T14 ? T8 : T1;
  assign T1 = T7 ? T5 : T2;
  assign T2 = T3 ? AcquireTracker_0_io_inner_release_ready : VoluntaryReleaseTracker_io_inner_release_ready;
  assign T3 = T4[1'h0:1'h0];
  assign T4 = release_idx;
  assign T5 = T6 ? AcquireTracker_2_io_inner_release_ready : AcquireTracker_1_io_inner_release_ready;
  assign T6 = T4[1'h0:1'h0];
  assign T7 = T4[1'h1:1'h1];
  assign T8 = T13 ? T11 : T9;
  assign T9 = T10 ? AcquireTracker_4_io_inner_release_ready : AcquireTracker_3_io_inner_release_ready;
  assign T10 = T4[1'h0:1'h0];
  assign T11 = T12 ? AcquireTracker_6_io_inner_release_ready : AcquireTracker_5_io_inner_release_ready;
  assign T12 = T4[1'h0:1'h0];
  assign T13 = T4[1'h1:1'h1];
  assign T14 = T4[2'h2:2'h2];
  assign io_inner_probe_bits_payload_p_type = probe_arb_io_out_bits_payload_p_type;
  assign io_inner_probe_bits_payload_master_xact_id = probe_arb_io_out_bits_payload_master_xact_id;
  assign io_inner_probe_bits_payload_addr = probe_arb_io_out_bits_payload_addr;
  assign io_inner_probe_bits_header_dst = probe_arb_io_out_bits_header_dst;
  assign io_inner_probe_bits_header_src = probe_arb_io_out_bits_header_src;
  assign io_inner_probe_valid = probe_arb_io_out_valid;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_grant_bits_payload_g_type = grant_arb_io_out_bits_payload_g_type;
  assign io_inner_grant_bits_payload_master_xact_id = grant_arb_io_out_bits_payload_master_xact_id;
  assign io_inner_grant_bits_payload_client_xact_id = grant_arb_io_out_bits_payload_client_xact_id;
  assign io_inner_grant_bits_payload_data = grant_arb_io_out_bits_payload_data;
  assign io_inner_grant_bits_header_dst = grant_arb_io_out_bits_header_dst;
  assign io_inner_grant_bits_header_src = grant_arb_io_out_bits_header_src;
  assign io_inner_grant_valid = grant_arb_io_out_valid;
  assign io_inner_acquire_ready = T15;
  assign T15 = T23 & T16;
  assign T16 = any_acquire_conflict ^ 1'h1;
  assign T23 = T24 | AcquireTracker_6_io_inner_acquire_ready;
  assign T24 = T25 | AcquireTracker_5_io_inner_acquire_ready;
  assign T25 = T26 | AcquireTracker_4_io_inner_acquire_ready;
  assign T26 = T27 | AcquireTracker_3_io_inner_acquire_ready;
  assign T27 = T28 | AcquireTracker_2_io_inner_acquire_ready;
  assign T28 = T29 | AcquireTracker_1_io_inner_acquire_ready;
  assign T29 = VoluntaryReleaseTracker_io_inner_acquire_ready | AcquireTracker_0_io_inner_acquire_ready;
  VoluntaryReleaseTracker VoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_0_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_0_ready ),
       .io_inner_grant_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_0_ready ),
       .io_inner_probe_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_header_src(  )
       //.io_inner_probe_bits_header_dst(  )
       //.io_inner_probe_bits_payload_addr(  )
       //.io_inner_probe_bits_payload_master_xact_id(  )
       //.io_inner_probe_bits_payload_p_type(  )
       .io_inner_release_ready( VoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( T55 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T54 ),
       .io_has_acquire_conflict( VoluntaryReleaseTracker_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_0 AcquireTracker_0(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_0_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_1_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_1_ready ),
       .io_inner_grant_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_1_ready ),
       .io_inner_probe_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_0_io_inner_release_ready ),
       .io_inner_release_valid( T52 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_0_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T51 ),
       .io_has_acquire_conflict( AcquireTracker_0_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_1 AcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_2_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_2_ready ),
       .io_inner_grant_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_2_ready ),
       .io_inner_probe_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( T49 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_1_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T48 ),
       .io_has_acquire_conflict( AcquireTracker_1_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_2 AcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_3_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_3_ready ),
       .io_inner_grant_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_3_ready ),
       .io_inner_probe_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( T46 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_2_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T45 ),
       .io_has_acquire_conflict( AcquireTracker_2_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_3 AcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_4_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_4_ready ),
       .io_inner_grant_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_4_ready ),
       .io_inner_probe_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( T43 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_3_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T42 ),
       .io_has_acquire_conflict( AcquireTracker_3_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_4 AcquireTracker_4(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_4_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_5_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_5_ready ),
       .io_inner_grant_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_4_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_5_ready ),
       .io_inner_probe_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_4_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_4_io_inner_release_ready ),
       .io_inner_release_valid( T40 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_4_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_4_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_4_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_4_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_5_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T39 ),
       .io_has_acquire_conflict( AcquireTracker_4_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_5 AcquireTracker_5(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_5_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_6_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_6_ready ),
       .io_inner_grant_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_5_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_6_ready ),
       .io_inner_probe_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_5_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_5_io_inner_release_ready ),
       .io_inner_release_valid( T37 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_5_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_5_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_5_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_5_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_6_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T36 ),
       .io_has_acquire_conflict( AcquireTracker_5_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_6 AcquireTracker_6(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_6_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_7_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_7_ready ),
       .io_inner_grant_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_6_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_7_ready ),
       .io_inner_probe_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_6_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_6_io_inner_release_ready ),
       .io_inner_release_valid( T34 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_6_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_6_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_6_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_6_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_7_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T32 ),
       .io_has_acquire_conflict( AcquireTracker_6_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  Arbiter_11 alloc_arb(
       .io_in_7_ready( alloc_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_acquire_ready ),
       //.io_in_7_bits(  )
       .io_in_6_ready( alloc_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_acquire_ready ),
       //.io_in_6_bits(  )
       .io_in_5_ready( alloc_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_acquire_ready ),
       //.io_in_5_bits(  )
       .io_in_4_ready( alloc_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_acquire_ready ),
       //.io_in_4_bits(  )
       .io_in_3_ready( alloc_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_acquire_ready ),
       //.io_in_3_bits(  )
       .io_in_2_ready( alloc_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_acquire_ready ),
       //.io_in_2_bits(  )
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_acquire_ready ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( T30 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_7_bits = {1{$random}};
    assign alloc_arb.io_in_6_bits = {1{$random}};
    assign alloc_arb.io_in_5_bits = {1{$random}};
    assign alloc_arb.io_in_4_bits = {1{$random}};
    assign alloc_arb.io_in_3_bits = {1{$random}};
    assign alloc_arb.io_in_2_bits = {1{$random}};
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  Arbiter_12 probe_arb(
       .io_in_7_ready( probe_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_in_7_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_in_7_bits_payload_master_xact_id( AcquireTracker_6_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_7_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_in_6_ready( probe_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_in_6_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_in_6_bits_payload_master_xact_id( AcquireTracker_5_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_6_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_in_5_ready( probe_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_in_5_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_in_5_bits_payload_master_xact_id( AcquireTracker_4_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_5_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_in_4_ready( probe_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_in_4_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_in_4_bits_payload_master_xact_id( AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_4_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_in_3_ready( probe_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_in_3_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_in_3_bits_payload_master_xact_id( AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_3_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_in_2_ready( probe_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_in_2_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_in_1_ready( probe_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_in_1_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_in_0_ready( probe_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       //.io_in_0_bits_payload_p_type(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( probe_arb_io_out_valid ),
       .io_out_bits_header_src( probe_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( probe_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( probe_arb_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( probe_arb_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( probe_arb_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign probe_arb.io_in_0_bits_header_src = {1{$random}};
    assign probe_arb.io_in_0_bits_header_dst = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_addr = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_master_xact_id = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_p_type = {1{$random}};
  `endif
  Arbiter_13 grant_arb(
       .io_in_7_ready( grant_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_in_7_bits_payload_data( AcquireTracker_6_io_inner_grant_bits_payload_data ),
       .io_in_7_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_master_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_7_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       .io_in_6_ready( grant_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_in_6_bits_payload_data( AcquireTracker_5_io_inner_grant_bits_payload_data ),
       .io_in_6_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_master_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_6_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       .io_in_5_ready( grant_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_in_5_bits_payload_data( AcquireTracker_4_io_inner_grant_bits_payload_data ),
       .io_in_5_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_master_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_5_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       .io_in_4_ready( grant_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_in_4_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_in_4_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_4_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       .io_in_3_ready( grant_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_in_3_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_in_3_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_3_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       .io_in_2_ready( grant_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_in_2_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       .io_in_1_ready( grant_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_in_1_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       .io_in_0_ready( grant_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_in_0_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_in_0_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( grant_arb_io_out_valid ),
       .io_out_bits_header_src( grant_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( grant_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_data( grant_arb_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( grant_arb_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( grant_arb_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( grant_arb_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  UncachedTileLinkIOArbiterThatPassesId outer_arb(.clk(clk), .reset(reset),
       .io_in_7_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_in_7_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       .io_in_7_acquire_bits_header_src( AcquireTracker_6_io_outer_acquire_bits_header_src ),
       //.io_in_7_acquire_bits_header_dst(  )
       .io_in_7_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_in_7_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_7_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_in_7_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_in_7_acquire_bits_payload_write_mask( AcquireTracker_6_io_outer_acquire_bits_payload_write_mask ),
       .io_in_7_acquire_bits_payload_subword_addr( AcquireTracker_6_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_7_acquire_bits_payload_atomic_opcode( AcquireTracker_6_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_7_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_in_7_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_in_7_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_in_7_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_in_7_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_in_7_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_in_7_grant_bits_payload_master_xact_id( outer_arb_io_in_7_grant_bits_payload_master_xact_id ),
       .io_in_7_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_in_7_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_in_7_finish_valid(  )
       //.io_in_7_finish_bits_header_src(  )
       //.io_in_7_finish_bits_header_dst(  )
       //.io_in_7_finish_bits_payload_master_xact_id(  )
       .io_in_6_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_in_6_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       .io_in_6_acquire_bits_header_src( AcquireTracker_5_io_outer_acquire_bits_header_src ),
       //.io_in_6_acquire_bits_header_dst(  )
       .io_in_6_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_in_6_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_6_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_in_6_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_in_6_acquire_bits_payload_write_mask( AcquireTracker_5_io_outer_acquire_bits_payload_write_mask ),
       .io_in_6_acquire_bits_payload_subword_addr( AcquireTracker_5_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_6_acquire_bits_payload_atomic_opcode( AcquireTracker_5_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_6_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_in_6_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_in_6_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_in_6_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_in_6_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_in_6_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_in_6_grant_bits_payload_master_xact_id( outer_arb_io_in_6_grant_bits_payload_master_xact_id ),
       .io_in_6_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_in_6_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_in_6_finish_valid(  )
       //.io_in_6_finish_bits_header_src(  )
       //.io_in_6_finish_bits_header_dst(  )
       //.io_in_6_finish_bits_payload_master_xact_id(  )
       .io_in_5_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_in_5_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       .io_in_5_acquire_bits_header_src( AcquireTracker_4_io_outer_acquire_bits_header_src ),
       //.io_in_5_acquire_bits_header_dst(  )
       .io_in_5_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_in_5_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_5_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_in_5_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_in_5_acquire_bits_payload_write_mask( AcquireTracker_4_io_outer_acquire_bits_payload_write_mask ),
       .io_in_5_acquire_bits_payload_subword_addr( AcquireTracker_4_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_5_acquire_bits_payload_atomic_opcode( AcquireTracker_4_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_5_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_in_5_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_in_5_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_in_5_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_in_5_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_in_5_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_in_5_grant_bits_payload_master_xact_id( outer_arb_io_in_5_grant_bits_payload_master_xact_id ),
       .io_in_5_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_in_5_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_in_5_finish_valid(  )
       //.io_in_5_finish_bits_header_src(  )
       //.io_in_5_finish_bits_header_dst(  )
       //.io_in_5_finish_bits_payload_master_xact_id(  )
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_in_4_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_in_4_acquire_bits_header_dst(  )
       .io_in_4_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_in_4_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_4_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_in_4_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_in_4_acquire_bits_payload_write_mask( AcquireTracker_3_io_outer_acquire_bits_payload_write_mask ),
       .io_in_4_acquire_bits_payload_subword_addr( AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_4_acquire_bits_payload_atomic_opcode( AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_4_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_in_4_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_in_4_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_in_4_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_in_4_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_in_4_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_in_4_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_in_4_finish_valid(  )
       //.io_in_4_finish_bits_header_src(  )
       //.io_in_4_finish_bits_header_dst(  )
       //.io_in_4_finish_bits_payload_master_xact_id(  )
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_in_3_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_in_3_acquire_bits_header_dst(  )
       .io_in_3_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_in_3_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_3_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_in_3_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_in_3_acquire_bits_payload_write_mask( AcquireTracker_2_io_outer_acquire_bits_payload_write_mask ),
       .io_in_3_acquire_bits_payload_subword_addr( AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_3_acquire_bits_payload_atomic_opcode( AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_3_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_in_3_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_in_3_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_in_3_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_in_3_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_in_3_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_in_3_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_in_3_finish_valid(  )
       //.io_in_3_finish_bits_header_src(  )
       //.io_in_3_finish_bits_header_dst(  )
       //.io_in_3_finish_bits_payload_master_xact_id(  )
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_in_2_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_in_2_acquire_bits_header_dst(  )
       .io_in_2_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_in_2_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_2_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_in_2_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_in_2_acquire_bits_payload_write_mask( AcquireTracker_1_io_outer_acquire_bits_payload_write_mask ),
       .io_in_2_acquire_bits_payload_subword_addr( AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_2_acquire_bits_payload_atomic_opcode( AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_2_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_in_2_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_in_2_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_in_2_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_in_2_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_in_2_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_in_2_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_in_2_finish_valid(  )
       //.io_in_2_finish_bits_header_src(  )
       //.io_in_2_finish_bits_header_dst(  )
       //.io_in_2_finish_bits_payload_master_xact_id(  )
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_in_1_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_write_mask( AcquireTracker_0_io_outer_acquire_bits_payload_write_mask ),
       .io_in_1_acquire_bits_payload_subword_addr( AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_1_acquire_bits_payload_atomic_opcode( AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_1_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_in_1_finish_valid(  )
       //.io_in_1_finish_bits_header_src(  )
       //.io_in_1_finish_bits_header_dst(  )
       //.io_in_1_finish_bits_payload_master_xact_id(  )
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_in_0_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_in_0_acquire_bits_header_dst(  )
       .io_in_0_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_write_mask( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask ),
       .io_in_0_acquire_bits_payload_subword_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_0_acquire_bits_payload_atomic_opcode( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_0_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_in_0_finish_valid(  )
       //.io_in_0_finish_bits_header_src(  )
       //.io_in_0_finish_bits_header_dst(  )
       //.io_in_0_finish_bits_payload_master_xact_id(  )
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( outer_arb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( outer_arb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( outer_arb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( outer_arb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( outer_arb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_a_type( outer_arb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_write_mask( outer_arb_io_out_acquire_bits_payload_write_mask ),
       .io_out_acquire_bits_payload_subword_addr( outer_arb_io_out_acquire_bits_payload_subword_addr ),
       .io_out_acquire_bits_payload_atomic_opcode( outer_arb_io_out_acquire_bits_payload_atomic_opcode ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_header_src( io_outer_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_outer_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_outer_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_outer_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_outer_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_g_type( io_outer_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_outer_finish_ready ),
       .io_out_finish_valid( outer_arb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( outer_arb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( outer_arb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( outer_arb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign outer_arb.io_in_7_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_valid = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_6_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_valid = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_5_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_valid = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_4_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_valid = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_3_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_valid = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_2_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_valid = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_1_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_valid = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_0_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_valid = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_payload_master_xact_id = {1{$random}};
  `endif
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire T10;
  wire[31:0] T11;
  reg [31:0] ram [1:0];
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[5:0] T15;
  wire[4:0] T16;
  wire[25:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_rw = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_addr, T15};
  assign T15 = {io_enq_bits_tag, io_enq_bits_rw};
  assign io_deq_bits_tag = T16;
  assign T16 = T11[3'h5:1'h1];
  assign io_deq_bits_addr = T17;
  assign T17 = T11[5'h1f:3'h6];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_13(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T16;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T17;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T18;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[127:0] T11;
  reg [127:0] ram [1:0];
  wire[127:0] T12;
  wire T13;
  wire empty;
  wire T14;
  wire T15;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T16 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T17 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T18 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign io_deq_valid = T13;
  assign T13 = empty ^ 1'h1;
  assign empty = ptr_match & T14;
  assign T14 = maybe_full ^ 1'h1;
  assign io_enq_ready = T15;
  assign T15 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits_data;
  end
endmodule

module MemIOUncachedTileLinkIOConverter(input clk, input reset,
    output io_uncached_acquire_ready,
    input  io_uncached_acquire_valid,
    input [1:0] io_uncached_acquire_bits_header_src,
    input [1:0] io_uncached_acquire_bits_header_dst,
    input [25:0] io_uncached_acquire_bits_payload_addr,
    input [1:0] io_uncached_acquire_bits_payload_client_xact_id,
    input [511:0] io_uncached_acquire_bits_payload_data,
    input [2:0] io_uncached_acquire_bits_payload_a_type,
    input [5:0] io_uncached_acquire_bits_payload_write_mask,
    input [2:0] io_uncached_acquire_bits_payload_subword_addr,
    input [3:0] io_uncached_acquire_bits_payload_atomic_opcode,
    input  io_uncached_grant_ready,
    output io_uncached_grant_valid,
    //output[1:0] io_uncached_grant_bits_header_src
    //output[1:0] io_uncached_grant_bits_header_dst
    output[511:0] io_uncached_grant_bits_payload_data,
    output[1:0] io_uncached_grant_bits_payload_client_xact_id,
    output[2:0] io_uncached_grant_bits_payload_master_xact_id,
    output[3:0] io_uncached_grant_bits_payload_g_type,
    //output io_uncached_finish_ready
    input  io_uncached_finish_valid,
    input [1:0] io_uncached_finish_bits_header_src,
    input [1:0] io_uncached_finish_bits_header_dst,
    input [2:0] io_uncached_finish_bits_payload_master_xact_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire[127:0] T56;
  reg [511:0] buf_out;
  wire[511:0] T57;
  wire[511:0] T58;
  wire T29;
  wire T30;
  reg  active_out;
  wire T53;
  wire T27;
  wire T28;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  reg [2:0] cnt_out;
  wire[2:0] T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T40;
  reg  has_data;
  wire T54;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  reg  cmd_sent_out;
  wire T55;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[511:0] T59;
  wire[383:0] T60;
  wire T38;
  wire T39;
  wire T61;
  wire T62;
  wire T63;
  wire[4:0] T64;
  reg [1:0] tag_out;
  wire[1:0] T65;
  reg [25:0] addr_out;
  wire[25:0] T66;
  wire T67;
  wire T68;
  wire T0;
  wire T1;
  reg [2:0] cnt_in;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  wire T5;
  reg  active_in;
  wire T51;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire[3:0] T14;
  wire[2:0] T15;
  wire[1:0] T16;
  wire[1:0] T52;
  reg [4:0] tag_in;
  wire[4:0] T17;
  wire[511:0] T18;
  reg [511:0] buf_in;
  wire[511:0] T19;
  wire[511:0] T20;
  wire[511:0] T21;
  wire[511:0] T22;
  wire[383:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire mem_cmd_q_io_enq_ready;
  wire mem_cmd_q_io_deq_valid;
  wire[25:0] mem_cmd_q_io_deq_bits_addr;
  wire[4:0] mem_cmd_q_io_deq_bits_tag;
  wire mem_cmd_q_io_deq_bits_rw;
  wire mem_data_q_io_enq_ready;
  wire mem_data_q_io_deq_valid;
  wire[127:0] mem_data_q_io_deq_bits_data;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    buf_out = {16{$random}};
    active_out = {1{$random}};
    cnt_out = {1{$random}};
    has_data = {1{$random}};
    cmd_sent_out = {1{$random}};
    tag_out = {1{$random}};
    addr_out = {1{$random}};
    cnt_in = {1{$random}};
    active_in = {1{$random}};
    tag_in = {1{$random}};
    buf_in = {16{$random}};
  end
`endif

  assign T56 = buf_out[7'h7f:1'h0];
  assign T57 = T38 ? T59 : T58;
  assign T58 = T29 ? io_uncached_acquire_bits_payload_data : buf_out;
  assign T29 = T30 & io_uncached_acquire_valid;
  assign T30 = active_out ^ 1'h1;
  assign T53 = reset ? 1'h0 : T27;
  assign T27 = T31 ? 1'h0 : T28;
  assign T28 = T29 ? 1'h1 : active_out;
  assign T31 = active_out & T32;
  assign T32 = cmd_sent_out & T33;
  assign T33 = T40 | T34;
  assign T34 = cnt_out == 3'h4;
  assign T35 = T38 ? T37 : T36;
  assign T36 = T29 ? 3'h0 : cnt_out;
  assign T37 = cnt_out + 3'h1;
  assign T40 = has_data ^ 1'h1;
  assign T54 = reset ? 1'h0 : T41;
  assign T41 = T29 ? T42 : has_data;
  assign T42 = T44 | T43;
  assign T43 = 3'h6 == io_uncached_acquire_bits_payload_a_type;
  assign T44 = T46 | T45;
  assign T45 = 3'h5 == io_uncached_acquire_bits_payload_a_type;
  assign T46 = 3'h3 == io_uncached_acquire_bits_payload_a_type;
  assign T55 = reset ? 1'h0 : T47;
  assign T47 = T49 ? 1'h1 : T48;
  assign T48 = T29 ? 1'h0 : cmd_sent_out;
  assign T49 = active_out & T50;
  assign T50 = mem_cmd_q_io_enq_ready & T67;
  assign T59 = {128'h0, T60};
  assign T60 = buf_out >> 8'h80;
  assign T38 = active_out & T39;
  assign T39 = mem_data_q_io_enq_ready & T61;
  assign T61 = T63 & T62;
  assign T62 = cnt_out < 3'h4;
  assign T63 = active_out & has_data;
  assign T64 = {3'h0, tag_out};
  assign T65 = T29 ? io_uncached_acquire_bits_payload_client_xact_id : tag_out;
  assign T66 = T29 ? io_uncached_acquire_bits_payload_addr : addr_out;
  assign T67 = active_out & T68;
  assign T68 = cmd_sent_out ^ 1'h1;
  assign io_mem_resp_ready = T0;
  assign T0 = T13 | T1;
  assign T1 = cnt_in < 3'h4;
  assign T2 = T11 ? T10 : T3;
  assign T3 = T4 ? 3'h1 : cnt_in;
  assign T4 = T5 & io_mem_resp_valid;
  assign T5 = active_in ^ 1'h1;
  assign T51 = reset ? 1'h0 : T6;
  assign T6 = T8 ? 1'h0 : T7;
  assign T7 = T4 ? 1'h1 : active_in;
  assign T8 = active_in & T9;
  assign T9 = io_uncached_grant_ready & io_uncached_grant_valid;
  assign T10 = cnt_in + 3'h1;
  assign T11 = active_in & T12;
  assign T12 = io_mem_resp_ready & io_mem_resp_valid;
  assign T13 = active_in ^ 1'h1;
  assign io_mem_req_data_bits_data = mem_data_q_io_deq_bits_data;
  assign io_mem_req_data_valid = mem_data_q_io_deq_valid;
  assign io_mem_req_cmd_bits_rw = mem_cmd_q_io_deq_bits_rw;
  assign io_mem_req_cmd_bits_tag = mem_cmd_q_io_deq_bits_tag;
  assign io_mem_req_cmd_bits_addr = mem_cmd_q_io_deq_bits_addr;
  assign io_mem_req_cmd_valid = mem_cmd_q_io_deq_valid;
  assign io_uncached_grant_bits_payload_g_type = T14;
  assign T14 = 4'h0;
  assign io_uncached_grant_bits_payload_master_xact_id = T15;
  assign T15 = 3'h0;
  assign io_uncached_grant_bits_payload_client_xact_id = T16;
  assign T16 = T52;
  assign T52 = tag_in[1'h1:1'h0];
  assign T17 = T4 ? io_mem_resp_bits_tag : tag_in;
  assign io_uncached_grant_bits_payload_data = T18;
  assign T18 = buf_in;
  assign T19 = T11 ? T22 : T20;
  assign T20 = T4 ? T21 : buf_in;
  assign T21 = io_mem_resp_bits_data << 9'h180;
  assign T22 = {io_mem_resp_bits_data, T23};
  assign T23 = buf_in[9'h1ff:8'h80];
  assign io_uncached_grant_valid = T24;
  assign T24 = active_in & T25;
  assign T25 = cnt_in == 3'h4;
  assign io_uncached_acquire_ready = T26;
  assign T26 = active_out ^ 1'h1;
  Queue_12 mem_cmd_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_cmd_q_io_enq_ready ),
       .io_enq_valid( T67 ),
       .io_enq_bits_addr( addr_out ),
       .io_enq_bits_tag( T64 ),
       .io_enq_bits_rw( has_data ),
       .io_deq_ready( io_mem_req_cmd_ready ),
       .io_deq_valid( mem_cmd_q_io_deq_valid ),
       .io_deq_bits_addr( mem_cmd_q_io_deq_bits_addr ),
       .io_deq_bits_tag( mem_cmd_q_io_deq_bits_tag ),
       .io_deq_bits_rw( mem_cmd_q_io_deq_bits_rw )
       //.io_count(  )
  );
  Queue_13 mem_data_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_data_q_io_enq_ready ),
       .io_enq_valid( T61 ),
       .io_enq_bits_data( T56 ),
       .io_deq_ready( io_mem_req_data_ready ),
       .io_deq_valid( mem_data_q_io_deq_valid ),
       .io_deq_bits_data( mem_data_q_io_deq_bits_data )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T38) begin
      buf_out <= T59;
    end else if(T29) begin
      buf_out <= io_uncached_acquire_bits_payload_data;
    end
    if(reset) begin
      active_out <= 1'h0;
    end else if(T31) begin
      active_out <= 1'h0;
    end else if(T29) begin
      active_out <= 1'h1;
    end
    if(T38) begin
      cnt_out <= T37;
    end else if(T29) begin
      cnt_out <= 3'h0;
    end
    if(reset) begin
      has_data <= 1'h0;
    end else if(T29) begin
      has_data <= T42;
    end
    if(reset) begin
      cmd_sent_out <= 1'h0;
    end else if(T49) begin
      cmd_sent_out <= 1'h1;
    end else if(T29) begin
      cmd_sent_out <= 1'h0;
    end
    if(T29) begin
      tag_out <= io_uncached_acquire_bits_payload_client_xact_id;
    end
    if(T29) begin
      addr_out <= io_uncached_acquire_bits_payload_addr;
    end
    if(T11) begin
      cnt_in <= T10;
    end else if(T4) begin
      cnt_in <= 3'h1;
    end
    if(reset) begin
      active_in <= 1'h0;
    end else if(T8) begin
      active_in <= 1'h0;
    end else if(T4) begin
      active_in <= 1'h1;
    end
    if(T4) begin
      tag_in <= io_mem_resp_bits_tag;
    end
    if(T11) begin
      buf_in <= T22;
    end else if(T4) begin
      buf_in <= T21;
    end
  end
endmodule

module HellaFlowQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
    //output[5:0] io_count
);

  wire[4:0] T0;
  wire[4:0] T1;
  wire[132:0] T2;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire atLeastTwo;
  wire T23;
  wire[4:0] T24;
  reg [4:0] deq_ptr;
  wire[4:0] T32;
  wire[4:0] T13;
  wire[4:0] T14;
  wire do_deq;
  wire T15;
  wire do_flow;
  wire T7;
  wire T16;
  reg [4:0] enq_ptr;
  wire[4:0] T33;
  wire[4:0] T9;
  wire[4:0] T10;
  wire do_enq;
  wire T6;
  wire T8;
  wire full;
  reg  maybe_full;
  wire T34;
  wire T25;
  wire T26;
  wire ptr_match;
  wire[4:0] T12;
  wire[4:0] T17;
  wire[132:0] T3;
  wire[132:0] T4;
  wire[132:0] T5;
  reg [4:0] ram_addr;
  wire[4:0] T11;
  wire empty;
  wire T27;
  wire[127:0] T28;
  wire[127:0] T29;
  wire T30;
  reg  ram_out_valid;
  wire T31;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    maybe_full = {1{$random}};
    ram_addr = {1{$random}};
    ram_out_valid = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = empty ? io_enq_bits_tag : T1;
  assign T1 = T2[3'h4:1'h0];
  assign T18 = io_deq_ready & T19;
  assign T19 = atLeastTwo | T20;
  assign T20 = T22 & T21;
  assign T21 = empty ^ 1'h1;
  assign T22 = io_deq_valid ^ 1'h1;
  assign atLeastTwo = full | T23;
  assign T23 = 5'h2 <= T24;
  assign T24 = enq_ptr - deq_ptr;
  assign T32 = reset ? 5'h0 : T13;
  assign T13 = do_deq ? T14 : deq_ptr;
  assign T14 = deq_ptr + 5'h1;
  assign do_deq = T16 & T15;
  assign T15 = do_flow ^ 1'h1;
  assign do_flow = T7;
  assign T7 = empty & io_deq_ready;
  assign T16 = io_deq_ready & io_deq_valid;
  assign T33 = reset ? 5'h0 : T9;
  assign T9 = do_enq ? T10 : enq_ptr;
  assign T10 = enq_ptr + 5'h1;
  assign do_enq = T8 & T6;
  assign T6 = do_flow ^ 1'h1;
  assign T8 = io_enq_ready & io_enq_valid;
  assign full = ptr_match & maybe_full;
  assign T34 = reset ? 1'h0 : T25;
  assign T25 = T26 ? do_enq : maybe_full;
  assign T26 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign T12 = io_deq_valid ? T17 : deq_ptr;
  assign T17 = deq_ptr + 5'h1;
  HellaFlowQueue_ram ram (
    .CLK(clk),
    .W0A(enq_ptr),
    .W0E(do_enq),
    .W0I(T4),
    .R1A(T12),
    .R1E(T18),
    .R1O(T2)
  );
  assign T4 = T5;
  assign T5 = {io_enq_bits_data, io_enq_bits_tag};
  assign T11 = T18 ? T12 : ram_addr;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_deq_bits_data = T28;
  assign T28 = empty ? io_enq_bits_data : T29;
  assign T29 = T2[8'h84:3'h5];
  assign io_deq_valid = T30;
  assign T30 = empty ? io_enq_valid : ram_out_valid;
  assign io_enq_ready = T31;
  assign T31 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      deq_ptr <= 5'h0;
    end else if(do_deq) begin
      deq_ptr <= T14;
    end
    if(reset) begin
      enq_ptr <= 5'h0;
    end else if(do_enq) begin
      enq_ptr <= T10;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T26) begin
      maybe_full <= do_enq;
    end
    if(T18) begin
      ram_addr <= T12;
    end
    ram_out_valid <= T18;
  end
endmodule

module Queue_15(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
);

  wire[4:0] T0;
  wire[132:0] T1;
  reg [132:0] ram [0:0];
  wire[132:0] T2;
  wire[132:0] T3;
  wire[132:0] T4;
  wire do_enq;
  wire[127:0] T5;
  wire T6;
  wire empty;
  reg  full;
  wire T11;
  wire T7;
  wire T8;
  wire do_deq;
  wire T9;
  wire T10;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {5{$random}};
    full = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = T1[3'h4:1'h0];
  assign T1 = ram[1'h0];
  assign T3 = T4;
  assign T4 = {io_enq_bits_data, io_enq_bits_tag};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_deq_bits_data = T5;
  assign T5 = T1[8'h84:3'h5];
  assign io_deq_valid = T6;
  assign T6 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign T11 = reset ? 1'h0 : T7;
  assign T7 = T8 ? do_enq : full;
  assign T8 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_enq_ready = T9;
  assign T9 = T10 | io_deq_ready;
  assign T10 = full ^ 1'h1;

  always @(posedge clk) begin
    if (do_enq)
      ram[1'h0] <= T3;
    if(reset) begin
      full <= 1'h0;
    end else if(T8) begin
      full <= do_enq;
    end
  end
endmodule

module HellaQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
    //output[5:0] io_count
);

  wire fq_io_enq_ready;
  wire fq_io_deq_valid;
  wire[127:0] fq_io_deq_bits_data;
  wire[4:0] fq_io_deq_bits_tag;
  wire Queue_16_io_enq_ready;
  wire Queue_16_io_deq_valid;
  wire[127:0] Queue_16_io_deq_bits_data;
  wire[4:0] Queue_16_io_deq_bits_tag;


  assign io_deq_bits_tag = Queue_16_io_deq_bits_tag;
  assign io_deq_bits_data = Queue_16_io_deq_bits_data;
  assign io_deq_valid = Queue_16_io_deq_valid;
  assign io_enq_ready = fq_io_enq_ready;
  HellaFlowQueue fq(.clk(clk), .reset(reset),
       .io_enq_ready( fq_io_enq_ready ),
       .io_enq_valid( io_enq_valid ),
       .io_enq_bits_data( io_enq_bits_data ),
       .io_enq_bits_tag( io_enq_bits_tag ),
       .io_deq_ready( Queue_16_io_enq_ready ),
       .io_deq_valid( fq_io_deq_valid ),
       .io_deq_bits_data( fq_io_deq_bits_data ),
       .io_deq_bits_tag( fq_io_deq_bits_tag )
       //.io_count(  )
  );
  Queue_15 Queue_16(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_16_io_enq_ready ),
       .io_enq_valid( fq_io_deq_valid ),
       .io_enq_bits_data( fq_io_deq_bits_data ),
       .io_enq_bits_tag( fq_io_deq_bits_tag ),
       .io_deq_ready( io_deq_ready ),
       .io_deq_valid( Queue_16_io_deq_valid ),
       .io_deq_bits_data( Queue_16_io_deq_bits_data ),
       .io_deq_bits_tag( Queue_16_io_deq_bits_tag )
  );
endmodule

module DRAMSideLLCNull(input clk, input reset,
    output io_cpu_req_cmd_ready,
    input  io_cpu_req_cmd_valid,
    input [25:0] io_cpu_req_cmd_bits_addr,
    input [4:0] io_cpu_req_cmd_bits_tag,
    input  io_cpu_req_cmd_bits_rw,
    output io_cpu_req_data_ready,
    input  io_cpu_req_data_valid,
    input [127:0] io_cpu_req_data_bits_data,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[127:0] io_cpu_resp_bits_data,
    output[4:0] io_cpu_resp_bits_tag,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire T0;
  wire cmdq_mask;
  wire watermark;
  reg [5:0] count;
  wire[5:0] T17;
  wire[5:0] T1;
  wire[5:0] T2;
  wire[5:0] T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire dec;
  wire T7;
  wire T8;
  wire T9;
  wire inc;
  wire T10;
  wire[5:0] T11;
  wire T12;
  wire T13;
  wire[5:0] T14;
  wire T15;
  wire T16;
  wire resp_dataq_io_deq_valid;
  wire[127:0] resp_dataq_io_deq_bits_data;
  wire[4:0] resp_dataq_io_deq_bits_tag;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    count = {1{$random}};
  end
`endif

  assign io_mem_req_data_bits_data = io_cpu_req_data_bits_data;
  assign io_mem_req_data_valid = io_cpu_req_data_valid;
  assign io_mem_req_cmd_bits_rw = io_cpu_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = io_cpu_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = io_cpu_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = T0;
  assign T0 = io_cpu_req_cmd_valid & cmdq_mask;
  assign cmdq_mask = io_cpu_req_cmd_bits_rw | watermark;
  assign watermark = 6'h4 <= count;
  assign T17 = reset ? 6'h20 : T1;
  assign T1 = T15 ? T14 : T2;
  assign T2 = T12 ? T11 : T3;
  assign T3 = T5 ? T4 : count;
  assign T4 = count + 6'h1;
  assign T5 = inc & T6;
  assign T6 = dec ^ 1'h1;
  assign dec = T7;
  assign T7 = T9 & T8;
  assign T8 = io_mem_req_cmd_bits_rw ^ 1'h1;
  assign T9 = io_mem_req_cmd_ready & io_mem_req_cmd_valid;
  assign inc = T10;
  assign T10 = io_cpu_resp_ready & resp_dataq_io_deq_valid;
  assign T11 = count - 6'h4;
  assign T12 = T13 & dec;
  assign T13 = inc ^ 1'h1;
  assign T14 = count - 6'h3;
  assign T15 = inc & dec;
  assign io_cpu_resp_bits_tag = resp_dataq_io_deq_bits_tag;
  assign io_cpu_resp_bits_data = resp_dataq_io_deq_bits_data;
  assign io_cpu_resp_valid = resp_dataq_io_deq_valid;
  assign io_cpu_req_data_ready = io_mem_req_data_ready;
  assign io_cpu_req_cmd_ready = T16;
  assign T16 = io_mem_req_cmd_ready & cmdq_mask;
  HellaQueue resp_dataq(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( io_mem_resp_valid ),
       .io_enq_bits_data( io_mem_resp_bits_data ),
       .io_enq_bits_tag( io_mem_resp_bits_tag ),
       .io_deq_ready( io_cpu_resp_ready ),
       .io_deq_valid( resp_dataq_io_deq_valid ),
       .io_deq_bits_data( resp_dataq_io_deq_bits_data ),
       .io_deq_bits_tag( resp_dataq_io_deq_bits_tag )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      count <= 6'h20;
    end else if(T15) begin
      count <= T14;
    end else if(T12) begin
      count <= T11;
    end else if(T5) begin
      count <= T4;
    end
  end
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] ram [1:0];
  wire[31:0] T2;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[5:0] T5;
  wire do_enq;
  reg  R6;
  wire T19;
  wire T7;
  wire T8;
  reg  R9;
  wire T20;
  wire T10;
  wire T11;
  wire do_deq;
  wire[4:0] T12;
  wire[25:0] T13;
  wire T14;
  wire empty;
  wire T15;
  reg  maybe_full;
  wire T21;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R6 = {1{$random}};
    R9 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_rw = T0;
  assign T0 = T1[1'h0:1'h0];
  assign T1 = ram[R9];
  assign T3 = T4;
  assign T4 = {io_enq_bits_addr, T5};
  assign T5 = {io_enq_bits_tag, io_enq_bits_rw};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R6;
  assign T8 = R6 + 1'h1;
  assign T20 = reset ? 1'h0 : T10;
  assign T10 = do_deq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_tag = T12;
  assign T12 = T1[3'h5:1'h1];
  assign io_deq_bits_addr = T13;
  assign T13 = T1[5'h1f:3'h6];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = ptr_match & T15;
  assign T15 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = R6 == R9;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T8;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_deq) begin
      R9 <= T11;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data
);

  wire[127:0] T0;
  wire[127:0] T1;
  reg [127:0] ram [3:0];
  wire[127:0] T2;
  wire do_enq;
  reg [1:0] R3;
  wire[1:0] T14;
  wire[1:0] T4;
  wire[1:0] T5;
  reg [1:0] R6;
  wire[1:0] T15;
  wire[1:0] T7;
  wire[1:0] T8;
  wire do_deq;
  wire T9;
  wire empty;
  wire T10;
  reg  maybe_full;
  wire T16;
  wire T11;
  wire T12;
  wire ptr_match;
  wire T13;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      ram[initvar] = {4{$random}};
    R3 = {1{$random}};
    R6 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[7'h7f:1'h0];
  assign T1 = ram[R6];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T14 = reset ? 2'h0 : T4;
  assign T4 = do_enq ? T5 : R3;
  assign T5 = R3 + 2'h1;
  assign T15 = reset ? 2'h0 : T7;
  assign T7 = do_deq ? T8 : R6;
  assign T8 = R6 + 2'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T9;
  assign T9 = empty ^ 1'h1;
  assign empty = ptr_match & T10;
  assign T10 = maybe_full ^ 1'h1;
  assign T16 = reset ? 1'h0 : T11;
  assign T11 = T12 ? do_enq : maybe_full;
  assign T12 = do_enq != do_deq;
  assign ptr_match = R3 == R6;
  assign io_enq_ready = T13;
  assign T13 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R3] <= io_enq_bits_data;
    if(reset) begin
      R3 <= 2'h0;
    end else if(do_enq) begin
      R3 <= T5;
    end
    if(reset) begin
      R6 <= 2'h0;
    end else if(do_deq) begin
      R6 <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T12) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module OuterMemorySystem(input clk, input reset,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [1:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input [2:0] io_tiles_0_acquire_bits_payload_a_type,
    input [5:0] io_tiles_0_acquire_bits_payload_write_mask,
    input [2:0] io_tiles_0_acquire_bits_payload_subword_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_atomic_opcode,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[1:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[2:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [2:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[2:0] io_tiles_0_probe_bits_payload_master_xact_id,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [1:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [2:0] io_tiles_0_release_bits_payload_master_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_acquire_ready,
    input  io_htif_acquire_valid,
    input [1:0] io_htif_acquire_bits_header_src,
    input [1:0] io_htif_acquire_bits_header_dst,
    input [25:0] io_htif_acquire_bits_payload_addr,
    input [1:0] io_htif_acquire_bits_payload_client_xact_id,
    input [511:0] io_htif_acquire_bits_payload_data,
    input [2:0] io_htif_acquire_bits_payload_a_type,
    input [5:0] io_htif_acquire_bits_payload_write_mask,
    input [2:0] io_htif_acquire_bits_payload_subword_addr,
    input [3:0] io_htif_acquire_bits_payload_atomic_opcode,
    input  io_htif_grant_ready,
    output io_htif_grant_valid,
    output[1:0] io_htif_grant_bits_header_src,
    output[1:0] io_htif_grant_bits_header_dst,
    output[511:0] io_htif_grant_bits_payload_data,
    output[1:0] io_htif_grant_bits_payload_client_xact_id,
    output[2:0] io_htif_grant_bits_payload_master_xact_id,
    output[3:0] io_htif_grant_bits_payload_g_type,
    output io_htif_finish_ready,
    input  io_htif_finish_valid,
    input [1:0] io_htif_finish_bits_header_src,
    input [1:0] io_htif_finish_bits_header_dst,
    input [2:0] io_htif_finish_bits_payload_master_xact_id,
    input  io_htif_probe_ready,
    output io_htif_probe_valid,
    output[1:0] io_htif_probe_bits_header_src,
    output[1:0] io_htif_probe_bits_header_dst,
    output[25:0] io_htif_probe_bits_payload_addr,
    output[2:0] io_htif_probe_bits_payload_master_xact_id,
    output[1:0] io_htif_probe_bits_payload_p_type,
    output io_htif_release_ready,
    input  io_htif_release_valid,
    input [1:0] io_htif_release_bits_header_src,
    input [1:0] io_htif_release_bits_header_dst,
    input [25:0] io_htif_release_bits_payload_addr,
    input [1:0] io_htif_release_bits_payload_client_xact_id,
    input [2:0] io_htif_release_bits_payload_master_xact_id,
    input [511:0] io_htif_release_bits_payload_data,
    input [2:0] io_htif_release_bits_payload_r_type,
    input  io_incoherent_1,
    input  io_incoherent_0,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire Queue_14_io_enq_ready;
  wire Queue_14_io_deq_valid;
  wire[25:0] Queue_14_io_deq_bits_addr;
  wire[4:0] Queue_14_io_deq_bits_tag;
  wire Queue_14_io_deq_bits_rw;
  wire Queue_15_io_enq_ready;
  wire Queue_15_io_deq_valid;
  wire[127:0] Queue_15_io_deq_bits_data;
  wire conv_io_uncached_acquire_ready;
  wire conv_io_uncached_grant_valid;
  wire[511:0] conv_io_uncached_grant_bits_payload_data;
  wire[1:0] conv_io_uncached_grant_bits_payload_client_xact_id;
  wire[2:0] conv_io_uncached_grant_bits_payload_master_xact_id;
  wire[3:0] conv_io_uncached_grant_bits_payload_g_type;
  wire conv_io_mem_req_cmd_valid;
  wire[25:0] conv_io_mem_req_cmd_bits_addr;
  wire[4:0] conv_io_mem_req_cmd_bits_tag;
  wire conv_io_mem_req_cmd_bits_rw;
  wire conv_io_mem_req_data_valid;
  wire[127:0] conv_io_mem_req_data_bits_data;
  wire conv_io_mem_resp_ready;
  wire net_io_clients_1_acquire_ready;
  wire net_io_clients_1_grant_valid;
  wire[1:0] net_io_clients_1_grant_bits_header_src;
  wire[1:0] net_io_clients_1_grant_bits_header_dst;
  wire[511:0] net_io_clients_1_grant_bits_payload_data;
  wire[1:0] net_io_clients_1_grant_bits_payload_client_xact_id;
  wire[2:0] net_io_clients_1_grant_bits_payload_master_xact_id;
  wire[3:0] net_io_clients_1_grant_bits_payload_g_type;
  wire net_io_clients_1_finish_ready;
  wire net_io_clients_1_probe_valid;
  wire[1:0] net_io_clients_1_probe_bits_header_src;
  wire[1:0] net_io_clients_1_probe_bits_header_dst;
  wire[25:0] net_io_clients_1_probe_bits_payload_addr;
  wire[2:0] net_io_clients_1_probe_bits_payload_master_xact_id;
  wire[1:0] net_io_clients_1_probe_bits_payload_p_type;
  wire net_io_clients_1_release_ready;
  wire net_io_clients_0_acquire_ready;
  wire net_io_clients_0_grant_valid;
  wire[1:0] net_io_clients_0_grant_bits_header_src;
  wire[1:0] net_io_clients_0_grant_bits_header_dst;
  wire[511:0] net_io_clients_0_grant_bits_payload_data;
  wire[1:0] net_io_clients_0_grant_bits_payload_client_xact_id;
  wire[2:0] net_io_clients_0_grant_bits_payload_master_xact_id;
  wire[3:0] net_io_clients_0_grant_bits_payload_g_type;
  wire net_io_clients_0_finish_ready;
  wire net_io_clients_0_probe_valid;
  wire[1:0] net_io_clients_0_probe_bits_header_src;
  wire[1:0] net_io_clients_0_probe_bits_header_dst;
  wire[25:0] net_io_clients_0_probe_bits_payload_addr;
  wire[2:0] net_io_clients_0_probe_bits_payload_master_xact_id;
  wire[1:0] net_io_clients_0_probe_bits_payload_p_type;
  wire net_io_clients_0_release_ready;
  wire net_io_masters_0_acquire_valid;
  wire[1:0] net_io_masters_0_acquire_bits_header_src;
  wire[1:0] net_io_masters_0_acquire_bits_header_dst;
  wire[25:0] net_io_masters_0_acquire_bits_payload_addr;
  wire[1:0] net_io_masters_0_acquire_bits_payload_client_xact_id;
  wire[511:0] net_io_masters_0_acquire_bits_payload_data;
  wire[2:0] net_io_masters_0_acquire_bits_payload_a_type;
  wire[5:0] net_io_masters_0_acquire_bits_payload_write_mask;
  wire[2:0] net_io_masters_0_acquire_bits_payload_subword_addr;
  wire[3:0] net_io_masters_0_acquire_bits_payload_atomic_opcode;
  wire net_io_masters_0_grant_ready;
  wire net_io_masters_0_finish_valid;
  wire[1:0] net_io_masters_0_finish_bits_header_src;
  wire[1:0] net_io_masters_0_finish_bits_header_dst;
  wire[2:0] net_io_masters_0_finish_bits_payload_master_xact_id;
  wire net_io_masters_0_probe_ready;
  wire net_io_masters_0_release_valid;
  wire[1:0] net_io_masters_0_release_bits_header_src;
  wire[1:0] net_io_masters_0_release_bits_header_dst;
  wire[25:0] net_io_masters_0_release_bits_payload_addr;
  wire[1:0] net_io_masters_0_release_bits_payload_client_xact_id;
  wire[2:0] net_io_masters_0_release_bits_payload_master_xact_id;
  wire[511:0] net_io_masters_0_release_bits_payload_data;
  wire[2:0] net_io_masters_0_release_bits_payload_r_type;
  wire L2CoherenceAgent_io_inner_acquire_ready;
  wire L2CoherenceAgent_io_inner_grant_valid;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_header_dst;
  wire[511:0] L2CoherenceAgent_io_inner_grant_bits_payload_data;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id;
  wire[2:0] L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id;
  wire[3:0] L2CoherenceAgent_io_inner_grant_bits_payload_g_type;
  wire L2CoherenceAgent_io_inner_finish_ready;
  wire L2CoherenceAgent_io_inner_probe_valid;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_header_dst;
  wire[25:0] L2CoherenceAgent_io_inner_probe_bits_payload_addr;
  wire[2:0] L2CoherenceAgent_io_inner_probe_bits_payload_master_xact_id;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_payload_p_type;
  wire L2CoherenceAgent_io_inner_release_ready;
  wire L2CoherenceAgent_io_outer_acquire_valid;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_header_dst;
  wire[25:0] L2CoherenceAgent_io_outer_acquire_bits_payload_addr;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id;
  wire[511:0] L2CoherenceAgent_io_outer_acquire_bits_payload_data;
  wire[2:0] L2CoherenceAgent_io_outer_acquire_bits_payload_a_type;
  wire[5:0] L2CoherenceAgent_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] L2CoherenceAgent_io_outer_acquire_bits_payload_subword_addr;
  wire[3:0] L2CoherenceAgent_io_outer_acquire_bits_payload_atomic_opcode;
  wire L2CoherenceAgent_io_outer_grant_ready;
  wire L2CoherenceAgent_io_outer_finish_valid;
  wire[1:0] L2CoherenceAgent_io_outer_finish_bits_header_src;
  wire[1:0] L2CoherenceAgent_io_outer_finish_bits_header_dst;
  wire[2:0] L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id;
  wire llc_io_cpu_req_cmd_ready;
  wire llc_io_cpu_req_data_ready;
  wire llc_io_cpu_resp_valid;
  wire[127:0] llc_io_cpu_resp_bits_data;
  wire[4:0] llc_io_cpu_resp_bits_tag;
  wire llc_io_mem_req_cmd_valid;
  wire[25:0] llc_io_mem_req_cmd_bits_addr;
  wire[4:0] llc_io_mem_req_cmd_bits_tag;
  wire llc_io_mem_req_cmd_bits_rw;
  wire llc_io_mem_req_data_valid;
  wire[127:0] llc_io_mem_req_data_bits_data;


  assign io_mem_req_data_bits_data = llc_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = llc_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = llc_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = llc_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = llc_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = llc_io_mem_req_cmd_valid;
  assign io_htif_release_ready = net_io_clients_1_release_ready;
  assign io_htif_probe_bits_payload_p_type = net_io_clients_1_probe_bits_payload_p_type;
  assign io_htif_probe_bits_payload_master_xact_id = net_io_clients_1_probe_bits_payload_master_xact_id;
  assign io_htif_probe_bits_payload_addr = net_io_clients_1_probe_bits_payload_addr;
  assign io_htif_probe_bits_header_dst = net_io_clients_1_probe_bits_header_dst;
  assign io_htif_probe_bits_header_src = net_io_clients_1_probe_bits_header_src;
  assign io_htif_probe_valid = net_io_clients_1_probe_valid;
  assign io_htif_finish_ready = net_io_clients_1_finish_ready;
  assign io_htif_grant_bits_payload_g_type = net_io_clients_1_grant_bits_payload_g_type;
  assign io_htif_grant_bits_payload_master_xact_id = net_io_clients_1_grant_bits_payload_master_xact_id;
  assign io_htif_grant_bits_payload_client_xact_id = net_io_clients_1_grant_bits_payload_client_xact_id;
  assign io_htif_grant_bits_payload_data = net_io_clients_1_grant_bits_payload_data;
  assign io_htif_grant_bits_header_dst = net_io_clients_1_grant_bits_header_dst;
  assign io_htif_grant_bits_header_src = net_io_clients_1_grant_bits_header_src;
  assign io_htif_grant_valid = net_io_clients_1_grant_valid;
  assign io_htif_acquire_ready = net_io_clients_1_acquire_ready;
  assign io_tiles_0_release_ready = net_io_clients_0_release_ready;
  assign io_tiles_0_probe_bits_payload_p_type = net_io_clients_0_probe_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_master_xact_id = net_io_clients_0_probe_bits_payload_master_xact_id;
  assign io_tiles_0_probe_bits_payload_addr = net_io_clients_0_probe_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = net_io_clients_0_probe_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = net_io_clients_0_probe_bits_header_src;
  assign io_tiles_0_probe_valid = net_io_clients_0_probe_valid;
  assign io_tiles_0_finish_ready = net_io_clients_0_finish_ready;
  assign io_tiles_0_grant_bits_payload_g_type = net_io_clients_0_grant_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_master_xact_id = net_io_clients_0_grant_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = net_io_clients_0_grant_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = net_io_clients_0_grant_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = net_io_clients_0_grant_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = net_io_clients_0_grant_bits_header_src;
  assign io_tiles_0_grant_valid = net_io_clients_0_grant_valid;
  assign io_tiles_0_acquire_ready = net_io_clients_0_acquire_ready;
  RocketChipCrossbarNetwork net(.clk(clk), .reset(reset),
       .io_clients_1_acquire_ready( net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( io_htif_acquire_valid ),
       .io_clients_1_acquire_bits_header_src( io_htif_acquire_bits_header_src ),
       .io_clients_1_acquire_bits_header_dst( io_htif_acquire_bits_header_dst ),
       .io_clients_1_acquire_bits_payload_addr( io_htif_acquire_bits_payload_addr ),
       .io_clients_1_acquire_bits_payload_client_xact_id( io_htif_acquire_bits_payload_client_xact_id ),
       .io_clients_1_acquire_bits_payload_data( io_htif_acquire_bits_payload_data ),
       .io_clients_1_acquire_bits_payload_a_type( io_htif_acquire_bits_payload_a_type ),
       .io_clients_1_acquire_bits_payload_write_mask( io_htif_acquire_bits_payload_write_mask ),
       .io_clients_1_acquire_bits_payload_subword_addr( io_htif_acquire_bits_payload_subword_addr ),
       .io_clients_1_acquire_bits_payload_atomic_opcode( io_htif_acquire_bits_payload_atomic_opcode ),
       .io_clients_1_grant_ready( io_htif_grant_ready ),
       .io_clients_1_grant_valid( net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_header_src( net_io_clients_1_grant_bits_header_src ),
       .io_clients_1_grant_bits_header_dst( net_io_clients_1_grant_bits_header_dst ),
       .io_clients_1_grant_bits_payload_data( net_io_clients_1_grant_bits_payload_data ),
       .io_clients_1_grant_bits_payload_client_xact_id( net_io_clients_1_grant_bits_payload_client_xact_id ),
       .io_clients_1_grant_bits_payload_master_xact_id( net_io_clients_1_grant_bits_payload_master_xact_id ),
       .io_clients_1_grant_bits_payload_g_type( net_io_clients_1_grant_bits_payload_g_type ),
       .io_clients_1_finish_ready( net_io_clients_1_finish_ready ),
       .io_clients_1_finish_valid( io_htif_finish_valid ),
       .io_clients_1_finish_bits_header_src( io_htif_finish_bits_header_src ),
       .io_clients_1_finish_bits_header_dst( io_htif_finish_bits_header_dst ),
       .io_clients_1_finish_bits_payload_master_xact_id( io_htif_finish_bits_payload_master_xact_id ),
       .io_clients_1_probe_ready( io_htif_probe_ready ),
       .io_clients_1_probe_valid( net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_header_src( net_io_clients_1_probe_bits_header_src ),
       .io_clients_1_probe_bits_header_dst( net_io_clients_1_probe_bits_header_dst ),
       .io_clients_1_probe_bits_payload_addr( net_io_clients_1_probe_bits_payload_addr ),
       .io_clients_1_probe_bits_payload_master_xact_id( net_io_clients_1_probe_bits_payload_master_xact_id ),
       .io_clients_1_probe_bits_payload_p_type( net_io_clients_1_probe_bits_payload_p_type ),
       .io_clients_1_release_ready( net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( io_htif_release_valid ),
       .io_clients_1_release_bits_header_src( io_htif_release_bits_header_src ),
       .io_clients_1_release_bits_header_dst( io_htif_release_bits_header_dst ),
       .io_clients_1_release_bits_payload_addr( io_htif_release_bits_payload_addr ),
       .io_clients_1_release_bits_payload_client_xact_id( io_htif_release_bits_payload_client_xact_id ),
       .io_clients_1_release_bits_payload_master_xact_id( io_htif_release_bits_payload_master_xact_id ),
       .io_clients_1_release_bits_payload_data( io_htif_release_bits_payload_data ),
       .io_clients_1_release_bits_payload_r_type( io_htif_release_bits_payload_r_type ),
       .io_clients_0_acquire_ready( net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_0_acquire_valid ),
       .io_clients_0_acquire_bits_header_src( io_tiles_0_acquire_bits_header_src ),
       .io_clients_0_acquire_bits_header_dst( io_tiles_0_acquire_bits_header_dst ),
       .io_clients_0_acquire_bits_payload_addr( io_tiles_0_acquire_bits_payload_addr ),
       .io_clients_0_acquire_bits_payload_client_xact_id( io_tiles_0_acquire_bits_payload_client_xact_id ),
       .io_clients_0_acquire_bits_payload_data( io_tiles_0_acquire_bits_payload_data ),
       .io_clients_0_acquire_bits_payload_a_type( io_tiles_0_acquire_bits_payload_a_type ),
       .io_clients_0_acquire_bits_payload_write_mask( io_tiles_0_acquire_bits_payload_write_mask ),
       .io_clients_0_acquire_bits_payload_subword_addr( io_tiles_0_acquire_bits_payload_subword_addr ),
       .io_clients_0_acquire_bits_payload_atomic_opcode( io_tiles_0_acquire_bits_payload_atomic_opcode ),
       .io_clients_0_grant_ready( io_tiles_0_grant_ready ),
       .io_clients_0_grant_valid( net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_header_src( net_io_clients_0_grant_bits_header_src ),
       .io_clients_0_grant_bits_header_dst( net_io_clients_0_grant_bits_header_dst ),
       .io_clients_0_grant_bits_payload_data( net_io_clients_0_grant_bits_payload_data ),
       .io_clients_0_grant_bits_payload_client_xact_id( net_io_clients_0_grant_bits_payload_client_xact_id ),
       .io_clients_0_grant_bits_payload_master_xact_id( net_io_clients_0_grant_bits_payload_master_xact_id ),
       .io_clients_0_grant_bits_payload_g_type( net_io_clients_0_grant_bits_payload_g_type ),
       .io_clients_0_finish_ready( net_io_clients_0_finish_ready ),
       .io_clients_0_finish_valid( io_tiles_0_finish_valid ),
       .io_clients_0_finish_bits_header_src( io_tiles_0_finish_bits_header_src ),
       .io_clients_0_finish_bits_header_dst( io_tiles_0_finish_bits_header_dst ),
       .io_clients_0_finish_bits_payload_master_xact_id( io_tiles_0_finish_bits_payload_master_xact_id ),
       .io_clients_0_probe_ready( io_tiles_0_probe_ready ),
       .io_clients_0_probe_valid( net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_header_src( net_io_clients_0_probe_bits_header_src ),
       .io_clients_0_probe_bits_header_dst( net_io_clients_0_probe_bits_header_dst ),
       .io_clients_0_probe_bits_payload_addr( net_io_clients_0_probe_bits_payload_addr ),
       .io_clients_0_probe_bits_payload_master_xact_id( net_io_clients_0_probe_bits_payload_master_xact_id ),
       .io_clients_0_probe_bits_payload_p_type( net_io_clients_0_probe_bits_payload_p_type ),
       .io_clients_0_release_ready( net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_0_release_valid ),
       .io_clients_0_release_bits_header_src( io_tiles_0_release_bits_header_src ),
       .io_clients_0_release_bits_header_dst( io_tiles_0_release_bits_header_dst ),
       .io_clients_0_release_bits_payload_addr( io_tiles_0_release_bits_payload_addr ),
       .io_clients_0_release_bits_payload_client_xact_id( io_tiles_0_release_bits_payload_client_xact_id ),
       .io_clients_0_release_bits_payload_master_xact_id( io_tiles_0_release_bits_payload_master_xact_id ),
       .io_clients_0_release_bits_payload_data( io_tiles_0_release_bits_payload_data ),
       .io_clients_0_release_bits_payload_r_type( io_tiles_0_release_bits_payload_r_type ),
       .io_masters_0_acquire_ready( L2CoherenceAgent_io_inner_acquire_ready ),
       .io_masters_0_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_masters_0_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_masters_0_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_masters_0_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_masters_0_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_masters_0_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_masters_0_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_masters_0_acquire_bits_payload_write_mask( net_io_masters_0_acquire_bits_payload_write_mask ),
       .io_masters_0_acquire_bits_payload_subword_addr( net_io_masters_0_acquire_bits_payload_subword_addr ),
       .io_masters_0_acquire_bits_payload_atomic_opcode( net_io_masters_0_acquire_bits_payload_atomic_opcode ),
       .io_masters_0_grant_ready( net_io_masters_0_grant_ready ),
       .io_masters_0_grant_valid( L2CoherenceAgent_io_inner_grant_valid ),
       .io_masters_0_grant_bits_header_src( L2CoherenceAgent_io_inner_grant_bits_header_src ),
       .io_masters_0_grant_bits_header_dst( L2CoherenceAgent_io_inner_grant_bits_header_dst ),
       .io_masters_0_grant_bits_payload_data( L2CoherenceAgent_io_inner_grant_bits_payload_data ),
       .io_masters_0_grant_bits_payload_client_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id ),
       .io_masters_0_grant_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id ),
       .io_masters_0_grant_bits_payload_g_type( L2CoherenceAgent_io_inner_grant_bits_payload_g_type ),
       .io_masters_0_finish_ready( L2CoherenceAgent_io_inner_finish_ready ),
       .io_masters_0_finish_valid( net_io_masters_0_finish_valid ),
       .io_masters_0_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_masters_0_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_masters_0_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_masters_0_probe_ready( net_io_masters_0_probe_ready ),
       .io_masters_0_probe_valid( L2CoherenceAgent_io_inner_probe_valid ),
       .io_masters_0_probe_bits_header_src( L2CoherenceAgent_io_inner_probe_bits_header_src ),
       .io_masters_0_probe_bits_header_dst( L2CoherenceAgent_io_inner_probe_bits_header_dst ),
       .io_masters_0_probe_bits_payload_addr( L2CoherenceAgent_io_inner_probe_bits_payload_addr ),
       .io_masters_0_probe_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_probe_bits_payload_master_xact_id ),
       .io_masters_0_probe_bits_payload_p_type( L2CoherenceAgent_io_inner_probe_bits_payload_p_type ),
       .io_masters_0_release_ready( L2CoherenceAgent_io_inner_release_ready ),
       .io_masters_0_release_valid( net_io_masters_0_release_valid ),
       .io_masters_0_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_masters_0_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_masters_0_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_masters_0_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_masters_0_release_bits_payload_master_xact_id( net_io_masters_0_release_bits_payload_master_xact_id ),
       .io_masters_0_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_masters_0_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type )
  );
  L2CoherenceAgent L2CoherenceAgent(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( L2CoherenceAgent_io_inner_acquire_ready ),
       .io_inner_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_inner_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( net_io_masters_0_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( net_io_masters_0_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( net_io_masters_0_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( net_io_masters_0_grant_ready ),
       .io_inner_grant_valid( L2CoherenceAgent_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( L2CoherenceAgent_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( L2CoherenceAgent_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( L2CoherenceAgent_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( L2CoherenceAgent_io_inner_grant_bits_payload_g_type ),
       .io_inner_finish_ready( L2CoherenceAgent_io_inner_finish_ready ),
       .io_inner_finish_valid( net_io_masters_0_finish_valid ),
       .io_inner_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( net_io_masters_0_probe_ready ),
       .io_inner_probe_valid( L2CoherenceAgent_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( L2CoherenceAgent_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( L2CoherenceAgent_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( L2CoherenceAgent_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( L2CoherenceAgent_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( L2CoherenceAgent_io_inner_release_ready ),
       .io_inner_release_valid( net_io_masters_0_release_valid ),
       .io_inner_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_inner_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( net_io_masters_0_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type ),
       .io_outer_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_outer_acquire_valid( L2CoherenceAgent_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( L2CoherenceAgent_io_outer_acquire_bits_header_src ),
       .io_outer_acquire_bits_header_dst( L2CoherenceAgent_io_outer_acquire_bits_header_dst ),
       .io_outer_acquire_bits_payload_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( L2CoherenceAgent_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( L2CoherenceAgent_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( L2CoherenceAgent_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( L2CoherenceAgent_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( L2CoherenceAgent_io_outer_grant_ready ),
       .io_outer_grant_valid( conv_io_uncached_grant_valid ),
       //.io_outer_grant_bits_header_src(  )
       //.io_outer_grant_bits_header_dst(  )
       .io_outer_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_outer_finish_ready(  )
       .io_outer_finish_valid( L2CoherenceAgent_io_outer_finish_valid ),
       .io_outer_finish_bits_header_src( L2CoherenceAgent_io_outer_finish_bits_header_src ),
       .io_outer_finish_bits_header_dst( L2CoherenceAgent_io_outer_finish_bits_header_dst ),
       .io_outer_finish_bits_payload_master_xact_id( L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id ),
       .io_incoherent_1( io_incoherent_1 ),
       .io_incoherent_0( io_incoherent_0 )
  );
  `ifndef SYNTHESIS
    assign L2CoherenceAgent.io_outer_grant_bits_header_src = {1{$random}};
    assign L2CoherenceAgent.io_outer_grant_bits_header_dst = {1{$random}};
    assign L2CoherenceAgent.io_outer_finish_ready = {1{$random}};
  `endif
  MemIOUncachedTileLinkIOConverter conv(.clk(clk), .reset(reset),
       .io_uncached_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_uncached_acquire_valid( L2CoherenceAgent_io_outer_acquire_valid ),
       .io_uncached_acquire_bits_header_src( L2CoherenceAgent_io_outer_acquire_bits_header_src ),
       .io_uncached_acquire_bits_header_dst( L2CoherenceAgent_io_outer_acquire_bits_header_dst ),
       .io_uncached_acquire_bits_payload_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_addr ),
       .io_uncached_acquire_bits_payload_client_xact_id( L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id ),
       .io_uncached_acquire_bits_payload_data( L2CoherenceAgent_io_outer_acquire_bits_payload_data ),
       .io_uncached_acquire_bits_payload_a_type( L2CoherenceAgent_io_outer_acquire_bits_payload_a_type ),
       .io_uncached_acquire_bits_payload_write_mask( L2CoherenceAgent_io_outer_acquire_bits_payload_write_mask ),
       .io_uncached_acquire_bits_payload_subword_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_subword_addr ),
       .io_uncached_acquire_bits_payload_atomic_opcode( L2CoherenceAgent_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_uncached_grant_ready( L2CoherenceAgent_io_outer_grant_ready ),
       .io_uncached_grant_valid( conv_io_uncached_grant_valid ),
       //.io_uncached_grant_bits_header_src(  )
       //.io_uncached_grant_bits_header_dst(  )
       .io_uncached_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_uncached_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_uncached_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_uncached_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_uncached_finish_ready(  )
       .io_uncached_finish_valid( L2CoherenceAgent_io_outer_finish_valid ),
       .io_uncached_finish_bits_header_src( L2CoherenceAgent_io_outer_finish_bits_header_src ),
       .io_uncached_finish_bits_header_dst( L2CoherenceAgent_io_outer_finish_bits_header_dst ),
       .io_uncached_finish_bits_payload_master_xact_id( L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id ),
       .io_mem_req_cmd_ready( Queue_14_io_enq_ready ),
       .io_mem_req_cmd_valid( conv_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( conv_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( conv_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( conv_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( Queue_15_io_enq_ready ),
       .io_mem_req_data_valid( conv_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( conv_io_mem_req_data_bits_data ),
       .io_mem_resp_ready( conv_io_mem_resp_ready ),
       .io_mem_resp_valid( llc_io_cpu_resp_valid ),
       .io_mem_resp_bits_data( llc_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_tag( llc_io_cpu_resp_bits_tag )
  );
  DRAMSideLLCNull llc(.clk(clk), .reset(reset),
       .io_cpu_req_cmd_ready( llc_io_cpu_req_cmd_ready ),
       .io_cpu_req_cmd_valid( Queue_14_io_deq_valid ),
       .io_cpu_req_cmd_bits_addr( Queue_14_io_deq_bits_addr ),
       .io_cpu_req_cmd_bits_tag( Queue_14_io_deq_bits_tag ),
       .io_cpu_req_cmd_bits_rw( Queue_14_io_deq_bits_rw ),
       .io_cpu_req_data_ready( llc_io_cpu_req_data_ready ),
       .io_cpu_req_data_valid( Queue_15_io_deq_valid ),
       .io_cpu_req_data_bits_data( Queue_15_io_deq_bits_data ),
       .io_cpu_resp_ready( conv_io_mem_resp_ready ),
       .io_cpu_resp_valid( llc_io_cpu_resp_valid ),
       .io_cpu_resp_bits_data( llc_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_tag( llc_io_cpu_resp_bits_tag ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( llc_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( llc_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( llc_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( llc_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( llc_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( llc_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
  );
  Queue_9 Queue_14(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_14_io_enq_ready ),
       .io_enq_valid( conv_io_mem_req_cmd_valid ),
       .io_enq_bits_addr( conv_io_mem_req_cmd_bits_addr ),
       .io_enq_bits_tag( conv_io_mem_req_cmd_bits_tag ),
       .io_enq_bits_rw( conv_io_mem_req_cmd_bits_rw ),
       .io_deq_ready( llc_io_cpu_req_cmd_ready ),
       .io_deq_valid( Queue_14_io_deq_valid ),
       .io_deq_bits_addr( Queue_14_io_deq_bits_addr ),
       .io_deq_bits_tag( Queue_14_io_deq_bits_tag ),
       .io_deq_bits_rw( Queue_14_io_deq_bits_rw )
  );
  Queue_10 Queue_15(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_15_io_enq_ready ),
       .io_enq_valid( conv_io_mem_req_data_valid ),
       .io_enq_bits_data( conv_io_mem_req_data_bits_data ),
       .io_deq_ready( llc_io_cpu_req_data_ready ),
       .io_deq_valid( Queue_15_io_deq_valid ),
       .io_deq_bits_data( Queue_15_io_deq_bits_data )
  );
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_a_type,
    input [5:0] io_enq_bits_payload_write_mask,
    input [2:0] io_enq_bits_payload_subword_addr,
    input [3:0] io_enq_bits_payload_atomic_opcode,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_a_type,
    output[5:0] io_deq_bits_payload_write_mask,
    output[2:0] io_deq_bits_payload_subword_addr,
    output[3:0] io_deq_bits_payload_atomic_opcode
);

  wire[3:0] T0;
  wire[559:0] T1;
  reg [559:0] ram [1:0];
  wire[559:0] T2;
  wire[559:0] T3;
  wire[559:0] T4;
  wire[527:0] T5;
  wire[12:0] T6;
  wire[6:0] T7;
  wire[514:0] T8;
  wire[31:0] T9;
  wire[27:0] T10;
  wire[3:0] T11;
  wire do_enq;
  reg  R12;
  wire T31;
  wire T13;
  wire T14;
  reg  R15;
  wire T32;
  wire T16;
  wire T17;
  wire do_deq;
  wire[2:0] T18;
  wire[5:0] T19;
  wire[2:0] T20;
  wire[511:0] T21;
  wire[1:0] T22;
  wire[25:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire empty;
  wire T27;
  reg  maybe_full;
  wire T33;
  wire T28;
  wire T29;
  wire ptr_match;
  wire T30;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {18{$random}};
    R12 = {1{$random}};
    R15 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_atomic_opcode = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = ram[R15];
  assign T3 = T4;
  assign T4 = {T9, T5};
  assign T5 = {T8, T6};
  assign T6 = {io_enq_bits_payload_write_mask, T7};
  assign T7 = {io_enq_bits_payload_subword_addr, io_enq_bits_payload_atomic_opcode};
  assign T8 = {io_enq_bits_payload_data, io_enq_bits_payload_a_type};
  assign T9 = {T11, T10};
  assign T10 = {io_enq_bits_payload_addr, io_enq_bits_payload_client_xact_id};
  assign T11 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T31 = reset ? 1'h0 : T13;
  assign T13 = do_enq ? T14 : R12;
  assign T14 = R12 + 1'h1;
  assign T32 = reset ? 1'h0 : T16;
  assign T16 = do_deq ? T17 : R15;
  assign T17 = R15 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_subword_addr = T18;
  assign T18 = T1[3'h6:3'h4];
  assign io_deq_bits_payload_write_mask = T19;
  assign T19 = T1[4'hc:3'h7];
  assign io_deq_bits_payload_a_type = T20;
  assign T20 = T1[4'hf:4'hd];
  assign io_deq_bits_payload_data = T21;
  assign T21 = T1[10'h20f:5'h10];
  assign io_deq_bits_payload_client_xact_id = T22;
  assign T22 = T1[10'h211:10'h210];
  assign io_deq_bits_payload_addr = T23;
  assign T23 = T1[10'h22b:10'h212];
  assign io_deq_bits_header_dst = T24;
  assign T24 = T1[10'h22d:10'h22c];
  assign io_deq_bits_header_src = T25;
  assign T25 = T1[10'h22f:10'h22e];
  assign io_deq_valid = T26;
  assign T26 = empty ^ 1'h1;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign T33 = reset ? 1'h0 : T28;
  assign T28 = T29 ? do_enq : maybe_full;
  assign T29 = do_enq != do_deq;
  assign ptr_match = R12 == R15;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R12] <= T3;
    if(reset) begin
      R12 <= 1'h0;
    end else if(do_enq) begin
      R12 <= T14;
    end
    if(reset) begin
      R15 <= 1'h0;
    end else if(do_deq) begin
      R15 <= T17;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T29) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_r_type
);

  wire[2:0] T0;
  wire[549:0] T1;
  reg [549:0] ram [1:0];
  wire[549:0] T2;
  wire[549:0] T3;
  wire[549:0] T4;
  wire[519:0] T5;
  wire[514:0] T6;
  wire[4:0] T7;
  wire[29:0] T8;
  wire[27:0] T9;
  wire do_enq;
  reg  R10;
  wire T27;
  wire T11;
  wire T12;
  reg  R13;
  wire T28;
  wire T14;
  wire T15;
  wire do_deq;
  wire[511:0] T16;
  wire[2:0] T17;
  wire[1:0] T18;
  wire[25:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire empty;
  wire T23;
  reg  maybe_full;
  wire T29;
  wire T24;
  wire T25;
  wire ptr_match;
  wire T26;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {18{$random}};
    R10 = {1{$random}};
    R13 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_r_type = T0;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = ram[R13];
  assign T3 = T4;
  assign T4 = {T8, T5};
  assign T5 = {T7, T6};
  assign T6 = {io_enq_bits_payload_data, io_enq_bits_payload_r_type};
  assign T7 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_master_xact_id};
  assign T8 = {io_enq_bits_header_src, T9};
  assign T9 = {io_enq_bits_header_dst, io_enq_bits_payload_addr};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T27 = reset ? 1'h0 : T11;
  assign T11 = do_enq ? T12 : R10;
  assign T12 = R10 + 1'h1;
  assign T28 = reset ? 1'h0 : T14;
  assign T14 = do_deq ? T15 : R13;
  assign T15 = R13 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_data = T16;
  assign T16 = T1[10'h202:2'h3];
  assign io_deq_bits_payload_master_xact_id = T17;
  assign T17 = T1[10'h205:10'h203];
  assign io_deq_bits_payload_client_xact_id = T18;
  assign T18 = T1[10'h207:10'h206];
  assign io_deq_bits_payload_addr = T19;
  assign T19 = T1[10'h221:10'h208];
  assign io_deq_bits_header_dst = T20;
  assign T20 = T1[10'h223:10'h222];
  assign io_deq_bits_header_src = T21;
  assign T21 = T1[10'h225:10'h224];
  assign io_deq_valid = T22;
  assign T22 = empty ^ 1'h1;
  assign empty = ptr_match & T23;
  assign T23 = maybe_full ^ 1'h1;
  assign T29 = reset ? 1'h0 : T24;
  assign T24 = T25 ? do_enq : maybe_full;
  assign T25 = do_enq != do_deq;
  assign ptr_match = R10 == R13;
  assign io_enq_ready = T26;
  assign T26 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R10] <= T3;
    if(reset) begin
      R10 <= 1'h0;
    end else if(do_enq) begin
      R10 <= T12;
    end
    if(reset) begin
      R13 <= 1'h0;
    end else if(do_deq) begin
      R13 <= T15;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T25) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_master_xact_id
);

  wire[2:0] T0;
  wire[6:0] T1;
  reg [6:0] ram [1:0];
  wire[6:0] T2;
  wire[6:0] T3;
  wire[6:0] T4;
  wire[4:0] T5;
  wire do_enq;
  reg  R6;
  wire T19;
  wire T7;
  wire T8;
  reg  R9;
  wire T20;
  wire T10;
  wire T11;
  wire do_deq;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire empty;
  wire T15;
  reg  maybe_full;
  wire T21;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R6 = {1{$random}};
    R9 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_master_xact_id = T0;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = ram[R9];
  assign T3 = T4;
  assign T4 = {io_enq_bits_header_src, T5};
  assign T5 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R6;
  assign T8 = R6 + 1'h1;
  assign T20 = reset ? 1'h0 : T10;
  assign T10 = do_deq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_header_dst = T12;
  assign T12 = T1[3'h4:2'h3];
  assign io_deq_bits_header_src = T13;
  assign T13 = T1[3'h6:3'h5];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = ptr_match & T15;
  assign T15 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = R6 == R9;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T8;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_deq) begin
      R9 <= T11;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [511:0] io_enq_bits_payload_data,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input [3:0] io_enq_bits_payload_g_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[511:0] io_deq_bits_payload_data,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output[3:0] io_deq_bits_payload_g_type
);

  wire[3:0] T0;
  wire[524:0] T1;
  reg [524:0] ram [0:0];
  wire[524:0] T2;
  wire[524:0] T3;
  wire[524:0] T4;
  wire[8:0] T5;
  wire[6:0] T6;
  wire[515:0] T7;
  wire[513:0] T8;
  wire do_enq;
  wire[2:0] T9;
  wire[1:0] T10;
  wire[511:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire empty;
  reg  full;
  wire T19;
  wire T15;
  wire T16;
  wire do_deq;
  wire T17;
  wire T18;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {17{$random}};
    full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_g_type = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = ram[1'h0];
  assign T3 = T4;
  assign T4 = {T7, T5};
  assign T5 = {io_enq_bits_payload_client_xact_id, T6};
  assign T6 = {io_enq_bits_payload_master_xact_id, io_enq_bits_payload_g_type};
  assign T7 = {io_enq_bits_header_src, T8};
  assign T8 = {io_enq_bits_header_dst, io_enq_bits_payload_data};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_deq_bits_payload_master_xact_id = T9;
  assign T9 = T1[3'h6:3'h4];
  assign io_deq_bits_payload_client_xact_id = T10;
  assign T10 = T1[4'h8:3'h7];
  assign io_deq_bits_payload_data = T11;
  assign T11 = T1[10'h208:4'h9];
  assign io_deq_bits_header_dst = T12;
  assign T12 = T1[10'h20a:10'h209];
  assign io_deq_bits_header_src = T13;
  assign T13 = T1[10'h20c:10'h20b];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign T19 = reset ? 1'h0 : T15;
  assign T15 = T16 ? do_enq : full;
  assign T16 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_enq_ready = T17;
  assign T17 = T18 | io_deq_ready;
  assign T18 = full ^ 1'h1;

  always @(posedge clk) begin
    if (do_enq)
      ram[1'h0] <= T3;
    if(reset) begin
      full <= 1'h0;
    end else if(T16) begin
      full <= do_enq;
    end
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output[1:0] io_deq_bits_payload_p_type
);

  wire[1:0] T0;
  wire[34:0] T1;
  reg [34:0] ram [1:0];
  wire[34:0] T2;
  wire[34:0] T3;
  wire[34:0] T4;
  wire[30:0] T5;
  wire[4:0] T6;
  wire[3:0] T7;
  wire do_enq;
  reg  R8;
  wire T23;
  wire T9;
  wire T10;
  reg  R11;
  wire T24;
  wire T12;
  wire T13;
  wire do_deq;
  wire[2:0] T14;
  wire[25:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire empty;
  wire T19;
  reg  maybe_full;
  wire T25;
  wire T20;
  wire T21;
  wire ptr_match;
  wire T22;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
    R8 = {1{$random}};
    R11 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_p_type = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = ram[R11];
  assign T3 = T4;
  assign T4 = {T7, T5};
  assign T5 = {io_enq_bits_payload_addr, T6};
  assign T6 = {io_enq_bits_payload_master_xact_id, io_enq_bits_payload_p_type};
  assign T7 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T23 = reset ? 1'h0 : T9;
  assign T9 = do_enq ? T10 : R8;
  assign T10 = R8 + 1'h1;
  assign T24 = reset ? 1'h0 : T12;
  assign T12 = do_deq ? T13 : R11;
  assign T13 = R11 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_master_xact_id = T14;
  assign T14 = T1[3'h4:2'h2];
  assign io_deq_bits_payload_addr = T15;
  assign T15 = T1[5'h1e:3'h5];
  assign io_deq_bits_header_dst = T16;
  assign T16 = T1[6'h20:5'h1f];
  assign io_deq_bits_header_src = T17;
  assign T17 = T1[6'h22:6'h21];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign T25 = reset ? 1'h0 : T20;
  assign T20 = T21 ? do_enq : maybe_full;
  assign T21 = do_enq != do_deq;
  assign ptr_match = R8 == R11;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R8] <= T3;
    if(reset) begin
      R8 <= 1'h0;
    end else if(do_enq) begin
      R8 <= T10;
    end
    if(reset) begin
      R11 <= 1'h0;
    end else if(do_deq) begin
      R11 <= T13;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T21) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Uncore(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [1:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input [2:0] io_tiles_0_acquire_bits_payload_a_type,
    input [5:0] io_tiles_0_acquire_bits_payload_write_mask,
    input [2:0] io_tiles_0_acquire_bits_payload_subword_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_atomic_opcode,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[1:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[2:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [2:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[2:0] io_tiles_0_probe_bits_payload_master_xact_id,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [1:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [2:0] io_tiles_0_release_bits_payload_master_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_0_reset,
    //output io_htif_0_id
    input  io_htif_0_pcr_req_ready,
    output io_htif_0_pcr_req_valid,
    output io_htif_0_pcr_req_bits_rw,
    output[4:0] io_htif_0_pcr_req_bits_addr,
    output[63:0] io_htif_0_pcr_req_bits_data,
    output io_htif_0_pcr_rep_ready,
    input  io_htif_0_pcr_rep_valid,
    input [63:0] io_htif_0_pcr_rep_bits,
    output io_htif_0_ipi_req_ready,
    input  io_htif_0_ipi_req_valid,
    input  io_htif_0_ipi_req_bits,
    input  io_htif_0_ipi_rep_ready,
    output io_htif_0_ipi_rep_valid,
    output io_htif_0_ipi_rep_bits,
    input  io_htif_0_debug_stats_pcr,
    input  io_incoherent_0
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire[2:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire[2:0] T7;
  wire[511:0] T8;
  wire[2:0] T9;
  wire[1:0] T10;
  wire[25:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire[3:0] T15;
  wire[2:0] T16;
  wire[5:0] T17;
  wire[2:0] T18;
  wire[511:0] T19;
  wire[1:0] T20;
  wire[25:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire[2:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire[2:0] T29;
  wire[511:0] T30;
  wire[2:0] T31;
  wire[1:0] T32;
  wire[25:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire T36;
  wire[3:0] T37;
  wire[2:0] T38;
  wire[5:0] T39;
  wire[2:0] T40;
  wire[511:0] T41;
  wire[1:0] T42;
  wire[25:0] T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T0;
  wire T1;
  wire T2;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_header_src;
  wire[1:0] Queue_4_io_deq_bits_header_dst;
  wire[25:0] Queue_4_io_deq_bits_payload_addr;
  wire[1:0] Queue_4_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_4_io_deq_bits_payload_data;
  wire[2:0] Queue_4_io_deq_bits_payload_a_type;
  wire[5:0] Queue_4_io_deq_bits_payload_write_mask;
  wire[2:0] Queue_4_io_deq_bits_payload_subword_addr;
  wire[3:0] Queue_4_io_deq_bits_payload_atomic_opcode;
  wire Queue_5_io_enq_ready;
  wire Queue_5_io_deq_valid;
  wire[1:0] Queue_5_io_deq_bits_header_src;
  wire[1:0] Queue_5_io_deq_bits_header_dst;
  wire[25:0] Queue_5_io_deq_bits_payload_addr;
  wire[1:0] Queue_5_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_5_io_deq_bits_payload_master_xact_id;
  wire[511:0] Queue_5_io_deq_bits_payload_data;
  wire[2:0] Queue_5_io_deq_bits_payload_r_type;
  wire Queue_6_io_enq_ready;
  wire Queue_6_io_deq_valid;
  wire[1:0] Queue_6_io_deq_bits_header_src;
  wire[1:0] Queue_6_io_deq_bits_header_dst;
  wire[2:0] Queue_6_io_deq_bits_payload_master_xact_id;
  wire Queue_7_io_enq_ready;
  wire Queue_7_io_deq_valid;
  wire[1:0] Queue_7_io_deq_bits_header_src;
  wire[1:0] Queue_7_io_deq_bits_header_dst;
  wire[511:0] Queue_7_io_deq_bits_payload_data;
  wire[1:0] Queue_7_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_7_io_deq_bits_payload_master_xact_id;
  wire[3:0] Queue_7_io_deq_bits_payload_g_type;
  wire Queue_8_io_enq_ready;
  wire Queue_8_io_deq_valid;
  wire[1:0] Queue_8_io_deq_bits_header_src;
  wire[1:0] Queue_8_io_deq_bits_header_dst;
  wire[25:0] Queue_8_io_deq_bits_payload_addr;
  wire[2:0] Queue_8_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_8_io_deq_bits_payload_p_type;
  wire Queue_9_io_enq_ready;
  wire Queue_9_io_deq_valid;
  wire[1:0] Queue_9_io_deq_bits_header_src;
  wire[1:0] Queue_9_io_deq_bits_header_dst;
  wire[25:0] Queue_9_io_deq_bits_payload_addr;
  wire[1:0] Queue_9_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_9_io_deq_bits_payload_data;
  wire[2:0] Queue_9_io_deq_bits_payload_a_type;
  wire[5:0] Queue_9_io_deq_bits_payload_write_mask;
  wire[2:0] Queue_9_io_deq_bits_payload_subword_addr;
  wire[3:0] Queue_9_io_deq_bits_payload_atomic_opcode;
  wire Queue_10_io_enq_ready;
  wire Queue_10_io_deq_valid;
  wire[1:0] Queue_10_io_deq_bits_header_src;
  wire[1:0] Queue_10_io_deq_bits_header_dst;
  wire[25:0] Queue_10_io_deq_bits_payload_addr;
  wire[1:0] Queue_10_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_10_io_deq_bits_payload_master_xact_id;
  wire[511:0] Queue_10_io_deq_bits_payload_data;
  wire[2:0] Queue_10_io_deq_bits_payload_r_type;
  wire Queue_11_io_enq_ready;
  wire Queue_11_io_deq_valid;
  wire[1:0] Queue_11_io_deq_bits_header_src;
  wire[1:0] Queue_11_io_deq_bits_header_dst;
  wire[2:0] Queue_11_io_deq_bits_payload_master_xact_id;
  wire Queue_12_io_enq_ready;
  wire Queue_12_io_deq_valid;
  wire[1:0] Queue_12_io_deq_bits_header_src;
  wire[1:0] Queue_12_io_deq_bits_header_dst;
  wire[511:0] Queue_12_io_deq_bits_payload_data;
  wire[1:0] Queue_12_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_12_io_deq_bits_payload_master_xact_id;
  wire[3:0] Queue_12_io_deq_bits_payload_g_type;
  wire Queue_13_io_enq_ready;
  wire Queue_13_io_deq_valid;
  wire[1:0] Queue_13_io_deq_bits_header_src;
  wire[1:0] Queue_13_io_deq_bits_header_dst;
  wire[25:0] Queue_13_io_deq_bits_payload_addr;
  wire[2:0] Queue_13_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_13_io_deq_bits_payload_p_type;
  wire htif_io_host_in_ready;
  wire htif_io_host_out_valid;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_debug_stats_pcr;
  wire htif_io_cpu_0_reset;
  wire htif_io_cpu_0_pcr_req_valid;
  wire htif_io_cpu_0_pcr_req_bits_rw;
  wire[4:0] htif_io_cpu_0_pcr_req_bits_addr;
  wire[63:0] htif_io_cpu_0_pcr_req_bits_data;
  wire htif_io_cpu_0_pcr_rep_ready;
  wire htif_io_cpu_0_ipi_req_ready;
  wire htif_io_cpu_0_ipi_rep_valid;
  wire htif_io_mem_acquire_valid;
  wire[25:0] htif_io_mem_acquire_bits_payload_addr;
  wire[1:0] htif_io_mem_acquire_bits_payload_client_xact_id;
  wire[511:0] htif_io_mem_acquire_bits_payload_data;
  wire[2:0] htif_io_mem_acquire_bits_payload_a_type;
  wire[5:0] htif_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] htif_io_mem_acquire_bits_payload_subword_addr;
  wire[3:0] htif_io_mem_acquire_bits_payload_atomic_opcode;
  wire htif_io_mem_grant_ready;
  wire htif_io_mem_finish_valid;
  wire[1:0] htif_io_mem_finish_bits_header_dst;
  wire[2:0] htif_io_mem_finish_bits_payload_master_xact_id;
  wire htif_io_mem_probe_ready;
  wire htif_io_mem_release_valid;
  wire[25:0] htif_io_mem_release_bits_payload_addr;
  wire[1:0] htif_io_mem_release_bits_payload_client_xact_id;
  wire[2:0] htif_io_mem_release_bits_payload_master_xact_id;
  wire[511:0] htif_io_mem_release_bits_payload_data;
  wire[2:0] htif_io_mem_release_bits_payload_r_type;
  wire outmemsys_io_tiles_0_acquire_ready;
  wire outmemsys_io_tiles_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_src;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_dst;
  wire[511:0] outmemsys_io_tiles_0_grant_bits_payload_data;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[2:0] outmemsys_io_tiles_0_grant_bits_payload_master_xact_id;
  wire[3:0] outmemsys_io_tiles_0_grant_bits_payload_g_type;
  wire outmemsys_io_tiles_0_finish_ready;
  wire outmemsys_io_tiles_0_probe_valid;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_src;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_dst;
  wire[25:0] outmemsys_io_tiles_0_probe_bits_payload_addr;
  wire[2:0] outmemsys_io_tiles_0_probe_bits_payload_master_xact_id;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_payload_p_type;
  wire outmemsys_io_tiles_0_release_ready;
  wire outmemsys_io_htif_acquire_ready;
  wire outmemsys_io_htif_grant_valid;
  wire[1:0] outmemsys_io_htif_grant_bits_header_src;
  wire[1:0] outmemsys_io_htif_grant_bits_header_dst;
  wire[511:0] outmemsys_io_htif_grant_bits_payload_data;
  wire[1:0] outmemsys_io_htif_grant_bits_payload_client_xact_id;
  wire[2:0] outmemsys_io_htif_grant_bits_payload_master_xact_id;
  wire[3:0] outmemsys_io_htif_grant_bits_payload_g_type;
  wire outmemsys_io_htif_finish_ready;
  wire outmemsys_io_htif_probe_valid;
  wire[1:0] outmemsys_io_htif_probe_bits_header_src;
  wire[1:0] outmemsys_io_htif_probe_bits_header_dst;
  wire[25:0] outmemsys_io_htif_probe_bits_payload_addr;
  wire[2:0] outmemsys_io_htif_probe_bits_payload_master_xact_id;
  wire[1:0] outmemsys_io_htif_probe_bits_payload_p_type;
  wire outmemsys_io_htif_release_ready;
  wire outmemsys_io_mem_req_cmd_valid;
  wire[25:0] outmemsys_io_mem_req_cmd_bits_addr;
  wire[4:0] outmemsys_io_mem_req_cmd_bits_tag;
  wire outmemsys_io_mem_req_cmd_bits_rw;
  wire outmemsys_io_mem_req_data_valid;
  wire[127:0] outmemsys_io_mem_req_data_bits_data;


  assign T3 = htif_io_mem_finish_bits_payload_master_xact_id;
  assign T4 = htif_io_mem_finish_bits_header_dst;
  assign T5 = 2'h1;
  assign T6 = htif_io_mem_finish_valid;
  assign T7 = htif_io_mem_release_bits_payload_r_type;
  assign T8 = htif_io_mem_release_bits_payload_data;
  assign T9 = htif_io_mem_release_bits_payload_master_xact_id;
  assign T10 = htif_io_mem_release_bits_payload_client_xact_id;
  assign T11 = htif_io_mem_release_bits_payload_addr;
  assign T12 = 2'h0;
  assign T13 = 2'h1;
  assign T14 = htif_io_mem_release_valid;
  assign T15 = htif_io_mem_acquire_bits_payload_atomic_opcode;
  assign T16 = htif_io_mem_acquire_bits_payload_subword_addr;
  assign T17 = htif_io_mem_acquire_bits_payload_write_mask;
  assign T18 = htif_io_mem_acquire_bits_payload_a_type;
  assign T19 = htif_io_mem_acquire_bits_payload_data;
  assign T20 = htif_io_mem_acquire_bits_payload_client_xact_id;
  assign T21 = htif_io_mem_acquire_bits_payload_addr;
  assign T22 = 2'h0;
  assign T23 = 2'h1;
  assign T24 = htif_io_mem_acquire_valid;
  assign T25 = io_tiles_0_finish_bits_payload_master_xact_id;
  assign T26 = io_tiles_0_finish_bits_header_dst;
  assign T27 = 2'h0;
  assign T28 = io_tiles_0_finish_valid;
  assign T29 = io_tiles_0_release_bits_payload_r_type;
  assign T30 = io_tiles_0_release_bits_payload_data;
  assign T31 = io_tiles_0_release_bits_payload_master_xact_id;
  assign T32 = io_tiles_0_release_bits_payload_client_xact_id;
  assign T33 = io_tiles_0_release_bits_payload_addr;
  assign T34 = 2'h0;
  assign T35 = 2'h0;
  assign T36 = io_tiles_0_release_valid;
  assign T37 = io_tiles_0_acquire_bits_payload_atomic_opcode;
  assign T38 = io_tiles_0_acquire_bits_payload_subword_addr;
  assign T39 = io_tiles_0_acquire_bits_payload_write_mask;
  assign T40 = io_tiles_0_acquire_bits_payload_a_type;
  assign T41 = io_tiles_0_acquire_bits_payload_data;
  assign T42 = io_tiles_0_acquire_bits_payload_client_xact_id;
  assign T43 = io_tiles_0_acquire_bits_payload_addr;
  assign T44 = 2'h0;
  assign T45 = 2'h0;
  assign T46 = io_tiles_0_acquire_valid;
  assign T47 = Queue_10_io_enq_ready;
  assign T48 = Queue_11_io_enq_ready;
  assign T49 = Queue_9_io_enq_ready;
  assign io_htif_0_ipi_rep_valid = htif_io_cpu_0_ipi_rep_valid;
  assign io_htif_0_ipi_req_ready = htif_io_cpu_0_ipi_req_ready;
  assign io_htif_0_pcr_rep_ready = htif_io_cpu_0_pcr_rep_ready;
  assign io_htif_0_pcr_req_bits_data = htif_io_cpu_0_pcr_req_bits_data;
  assign io_htif_0_pcr_req_bits_addr = htif_io_cpu_0_pcr_req_bits_addr;
  assign io_htif_0_pcr_req_bits_rw = htif_io_cpu_0_pcr_req_bits_rw;
  assign io_htif_0_pcr_req_valid = htif_io_cpu_0_pcr_req_valid;
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign io_tiles_0_release_ready = T0;
  assign T0 = Queue_5_io_enq_ready;
  assign io_tiles_0_probe_bits_payload_p_type = Queue_8_io_deq_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_master_xact_id = Queue_8_io_deq_bits_payload_master_xact_id;
  assign io_tiles_0_probe_bits_payload_addr = Queue_8_io_deq_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = Queue_8_io_deq_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = Queue_8_io_deq_bits_header_src;
  assign io_tiles_0_probe_valid = Queue_8_io_deq_valid;
  assign io_tiles_0_finish_ready = T1;
  assign T1 = Queue_6_io_enq_ready;
  assign io_tiles_0_grant_bits_payload_g_type = Queue_7_io_deq_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_master_xact_id = Queue_7_io_deq_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = Queue_7_io_deq_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = Queue_7_io_deq_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = Queue_7_io_deq_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = Queue_7_io_deq_bits_header_src;
  assign io_tiles_0_grant_valid = Queue_7_io_deq_valid;
  assign io_tiles_0_acquire_ready = T2;
  assign T2 = Queue_4_io_enq_ready;
  assign io_mem_req_data_bits_data = outmemsys_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = outmemsys_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = outmemsys_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = outmemsys_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = outmemsys_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = outmemsys_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = htif_io_host_debug_stats_pcr;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_in_ready = htif_io_host_in_ready;
  HTIF htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       .io_host_debug_stats_pcr( htif_io_host_debug_stats_pcr ),
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       //.io_cpu_0_id(  )
       .io_cpu_0_pcr_req_ready( io_htif_0_pcr_req_ready ),
       .io_cpu_0_pcr_req_valid( htif_io_cpu_0_pcr_req_valid ),
       .io_cpu_0_pcr_req_bits_rw( htif_io_cpu_0_pcr_req_bits_rw ),
       .io_cpu_0_pcr_req_bits_addr( htif_io_cpu_0_pcr_req_bits_addr ),
       .io_cpu_0_pcr_req_bits_data( htif_io_cpu_0_pcr_req_bits_data ),
       .io_cpu_0_pcr_rep_ready( htif_io_cpu_0_pcr_rep_ready ),
       .io_cpu_0_pcr_rep_valid( io_htif_0_pcr_rep_valid ),
       .io_cpu_0_pcr_rep_bits( io_htif_0_pcr_rep_bits ),
       .io_cpu_0_ipi_req_ready( htif_io_cpu_0_ipi_req_ready ),
       .io_cpu_0_ipi_req_valid( io_htif_0_ipi_req_valid ),
       .io_cpu_0_ipi_req_bits( io_htif_0_ipi_req_bits ),
       .io_cpu_0_ipi_rep_ready( io_htif_0_ipi_rep_ready ),
       .io_cpu_0_ipi_rep_valid( htif_io_cpu_0_ipi_rep_valid ),
       //.io_cpu_0_ipi_rep_bits(  )
       .io_cpu_0_debug_stats_pcr( io_htif_0_debug_stats_pcr ),
       .io_mem_acquire_ready( T49 ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( htif_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( htif_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( htif_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( htif_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( htif_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( htif_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( htif_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( Queue_12_io_deq_valid ),
       .io_mem_grant_bits_header_src( Queue_12_io_deq_bits_header_src ),
       .io_mem_grant_bits_header_dst( Queue_12_io_deq_bits_header_dst ),
       .io_mem_grant_bits_payload_data( Queue_12_io_deq_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( Queue_12_io_deq_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( Queue_12_io_deq_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( Queue_12_io_deq_bits_payload_g_type ),
       .io_mem_finish_ready( T48 ),
       .io_mem_finish_valid( htif_io_mem_finish_valid ),
       //.io_mem_finish_bits_header_src(  )
       .io_mem_finish_bits_header_dst( htif_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( htif_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( htif_io_mem_probe_ready ),
       .io_mem_probe_valid( Queue_13_io_deq_valid ),
       .io_mem_probe_bits_header_src( Queue_13_io_deq_bits_header_src ),
       .io_mem_probe_bits_header_dst( Queue_13_io_deq_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( Queue_13_io_deq_bits_payload_addr ),
       .io_mem_probe_bits_payload_master_xact_id( Queue_13_io_deq_bits_payload_master_xact_id ),
       .io_mem_probe_bits_payload_p_type( Queue_13_io_deq_bits_payload_p_type ),
       .io_mem_release_ready( T47 ),
       .io_mem_release_valid( htif_io_mem_release_valid ),
       //.io_mem_release_bits_header_src(  )
       //.io_mem_release_bits_header_dst(  )
       .io_mem_release_bits_payload_addr( htif_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( htif_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_master_xact_id( htif_io_mem_release_bits_payload_master_xact_id ),
       .io_mem_release_bits_payload_data( htif_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( htif_io_mem_release_bits_payload_r_type )
       //.io_scr_rdata_63(  )
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       //.io_scr_rdata_2(  )
       //.io_scr_rdata_1(  )
       //.io_scr_rdata_0(  )
       //.io_scr_wen(  )
       //.io_scr_waddr(  )
       //.io_scr_wdata(  )
  );
  `ifndef SYNTHESIS
    assign htif.io_mem_release_bits_payload_addr = {1{$random}};
    assign htif.io_mem_release_bits_payload_client_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_master_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_data = {16{$random}};
    assign htif.io_mem_release_bits_payload_r_type = {1{$random}};
    assign htif.io_scr_rdata_63 = {2{$random}};
    assign htif.io_scr_rdata_62 = {2{$random}};
    assign htif.io_scr_rdata_61 = {2{$random}};
    assign htif.io_scr_rdata_60 = {2{$random}};
    assign htif.io_scr_rdata_59 = {2{$random}};
    assign htif.io_scr_rdata_58 = {2{$random}};
    assign htif.io_scr_rdata_57 = {2{$random}};
    assign htif.io_scr_rdata_56 = {2{$random}};
    assign htif.io_scr_rdata_55 = {2{$random}};
    assign htif.io_scr_rdata_54 = {2{$random}};
    assign htif.io_scr_rdata_53 = {2{$random}};
    assign htif.io_scr_rdata_52 = {2{$random}};
    assign htif.io_scr_rdata_51 = {2{$random}};
    assign htif.io_scr_rdata_50 = {2{$random}};
    assign htif.io_scr_rdata_49 = {2{$random}};
    assign htif.io_scr_rdata_48 = {2{$random}};
    assign htif.io_scr_rdata_47 = {2{$random}};
    assign htif.io_scr_rdata_46 = {2{$random}};
    assign htif.io_scr_rdata_45 = {2{$random}};
    assign htif.io_scr_rdata_44 = {2{$random}};
    assign htif.io_scr_rdata_43 = {2{$random}};
    assign htif.io_scr_rdata_42 = {2{$random}};
    assign htif.io_scr_rdata_41 = {2{$random}};
    assign htif.io_scr_rdata_40 = {2{$random}};
    assign htif.io_scr_rdata_39 = {2{$random}};
    assign htif.io_scr_rdata_38 = {2{$random}};
    assign htif.io_scr_rdata_37 = {2{$random}};
    assign htif.io_scr_rdata_36 = {2{$random}};
    assign htif.io_scr_rdata_35 = {2{$random}};
    assign htif.io_scr_rdata_34 = {2{$random}};
    assign htif.io_scr_rdata_33 = {2{$random}};
    assign htif.io_scr_rdata_32 = {2{$random}};
    assign htif.io_scr_rdata_31 = {2{$random}};
    assign htif.io_scr_rdata_30 = {2{$random}};
    assign htif.io_scr_rdata_29 = {2{$random}};
    assign htif.io_scr_rdata_28 = {2{$random}};
    assign htif.io_scr_rdata_27 = {2{$random}};
    assign htif.io_scr_rdata_26 = {2{$random}};
    assign htif.io_scr_rdata_25 = {2{$random}};
    assign htif.io_scr_rdata_24 = {2{$random}};
    assign htif.io_scr_rdata_23 = {2{$random}};
    assign htif.io_scr_rdata_22 = {2{$random}};
    assign htif.io_scr_rdata_21 = {2{$random}};
    assign htif.io_scr_rdata_20 = {2{$random}};
    assign htif.io_scr_rdata_19 = {2{$random}};
    assign htif.io_scr_rdata_18 = {2{$random}};
    assign htif.io_scr_rdata_17 = {2{$random}};
    assign htif.io_scr_rdata_16 = {2{$random}};
    assign htif.io_scr_rdata_15 = {2{$random}};
    assign htif.io_scr_rdata_14 = {2{$random}};
    assign htif.io_scr_rdata_13 = {2{$random}};
    assign htif.io_scr_rdata_12 = {2{$random}};
    assign htif.io_scr_rdata_11 = {2{$random}};
    assign htif.io_scr_rdata_10 = {2{$random}};
    assign htif.io_scr_rdata_9 = {2{$random}};
    assign htif.io_scr_rdata_8 = {2{$random}};
    assign htif.io_scr_rdata_7 = {2{$random}};
    assign htif.io_scr_rdata_6 = {2{$random}};
    assign htif.io_scr_rdata_5 = {2{$random}};
    assign htif.io_scr_rdata_4 = {2{$random}};
    assign htif.io_scr_rdata_3 = {2{$random}};
    assign htif.io_scr_rdata_2 = {2{$random}};
  `endif
  OuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_0_acquire_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( Queue_4_io_deq_valid ),
       .io_tiles_0_acquire_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( Queue_4_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( Queue_4_io_deq_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_a_type( Queue_4_io_deq_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_write_mask( Queue_4_io_deq_bits_payload_write_mask ),
       .io_tiles_0_acquire_bits_payload_subword_addr( Queue_4_io_deq_bits_payload_subword_addr ),
       .io_tiles_0_acquire_bits_payload_atomic_opcode( Queue_4_io_deq_bits_payload_atomic_opcode ),
       .io_tiles_0_grant_ready( Queue_7_io_enq_ready ),
       .io_tiles_0_grant_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( Queue_6_io_deq_valid ),
       .io_tiles_0_finish_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( Queue_8_io_enq_ready ),
       .io_tiles_0_probe_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_master_xact_id( outmemsys_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tiles_0_probe_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( outmemsys_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( Queue_5_io_deq_valid ),
       .io_tiles_0_release_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_master_xact_id( Queue_5_io_deq_bits_payload_master_xact_id ),
       .io_tiles_0_release_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( Queue_5_io_deq_bits_payload_r_type ),
       .io_htif_acquire_ready( outmemsys_io_htif_acquire_ready ),
       .io_htif_acquire_valid( Queue_9_io_deq_valid ),
       .io_htif_acquire_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_htif_acquire_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_htif_acquire_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_htif_acquire_bits_payload_client_xact_id( Queue_9_io_deq_bits_payload_client_xact_id ),
       .io_htif_acquire_bits_payload_data( Queue_9_io_deq_bits_payload_data ),
       .io_htif_acquire_bits_payload_a_type( Queue_9_io_deq_bits_payload_a_type ),
       .io_htif_acquire_bits_payload_write_mask( Queue_9_io_deq_bits_payload_write_mask ),
       .io_htif_acquire_bits_payload_subword_addr( Queue_9_io_deq_bits_payload_subword_addr ),
       .io_htif_acquire_bits_payload_atomic_opcode( Queue_9_io_deq_bits_payload_atomic_opcode ),
       .io_htif_grant_ready( Queue_12_io_enq_ready ),
       .io_htif_grant_valid( outmemsys_io_htif_grant_valid ),
       .io_htif_grant_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_htif_grant_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_htif_grant_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_htif_grant_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_htif_grant_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_htif_grant_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_htif_finish_ready( outmemsys_io_htif_finish_ready ),
       .io_htif_finish_valid( Queue_11_io_deq_valid ),
       .io_htif_finish_bits_header_src( Queue_11_io_deq_bits_header_src ),
       .io_htif_finish_bits_header_dst( Queue_11_io_deq_bits_header_dst ),
       .io_htif_finish_bits_payload_master_xact_id( Queue_11_io_deq_bits_payload_master_xact_id ),
       .io_htif_probe_ready( Queue_13_io_enq_ready ),
       .io_htif_probe_valid( outmemsys_io_htif_probe_valid ),
       .io_htif_probe_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_htif_probe_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_htif_probe_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_htif_probe_bits_payload_master_xact_id( outmemsys_io_htif_probe_bits_payload_master_xact_id ),
       .io_htif_probe_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_htif_release_ready( outmemsys_io_htif_release_ready ),
       .io_htif_release_valid( Queue_10_io_deq_valid ),
       .io_htif_release_bits_header_src( Queue_10_io_deq_bits_header_src ),
       .io_htif_release_bits_header_dst( Queue_10_io_deq_bits_header_dst ),
       .io_htif_release_bits_payload_addr( Queue_10_io_deq_bits_payload_addr ),
       .io_htif_release_bits_payload_client_xact_id( Queue_10_io_deq_bits_payload_client_xact_id ),
       .io_htif_release_bits_payload_master_xact_id( Queue_10_io_deq_bits_payload_master_xact_id ),
       .io_htif_release_bits_payload_data( Queue_10_io_deq_bits_payload_data ),
       .io_htif_release_bits_payload_r_type( Queue_10_io_deq_bits_payload_r_type ),
       .io_incoherent_1( 1'h1 ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( outmemsys_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( outmemsys_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( outmemsys_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( outmemsys_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( outmemsys_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( outmemsys_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
  Queue_3 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( T46 ),
       .io_enq_bits_header_src( T45 ),
       .io_enq_bits_header_dst( T44 ),
       .io_enq_bits_payload_addr( T43 ),
       .io_enq_bits_payload_client_xact_id( T42 ),
       .io_enq_bits_payload_data( T41 ),
       .io_enq_bits_payload_a_type( T40 ),
       .io_enq_bits_payload_write_mask( T39 ),
       .io_enq_bits_payload_subword_addr( T38 ),
       .io_enq_bits_payload_atomic_opcode( T37 ),
       .io_deq_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_4_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_4_io_deq_bits_payload_data ),
       .io_deq_bits_payload_a_type( Queue_4_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_write_mask( Queue_4_io_deq_bits_payload_write_mask ),
       .io_deq_bits_payload_subword_addr( Queue_4_io_deq_bits_payload_subword_addr ),
       .io_deq_bits_payload_atomic_opcode( Queue_4_io_deq_bits_payload_atomic_opcode )
  );
  Queue_4 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( T36 ),
       .io_enq_bits_header_src( T35 ),
       .io_enq_bits_header_dst( T34 ),
       .io_enq_bits_payload_addr( T33 ),
       .io_enq_bits_payload_client_xact_id( T32 ),
       .io_enq_bits_payload_master_xact_id( T31 ),
       .io_enq_bits_payload_data( T30 ),
       .io_enq_bits_payload_r_type( T29 ),
       .io_deq_ready( outmemsys_io_tiles_0_release_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_5_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_5_io_deq_bits_payload_r_type )
  );
  Queue_5 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( T28 ),
       .io_enq_bits_header_src( T27 ),
       .io_enq_bits_header_dst( T26 ),
       .io_enq_bits_payload_master_xact_id( T25 ),
       .io_deq_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id )
  );
  Queue_6 Queue_7(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_7_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_deq_ready( io_tiles_0_grant_ready ),
       .io_deq_valid( Queue_7_io_deq_valid ),
       .io_deq_bits_header_src( Queue_7_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_7_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_7_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_7_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_7_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_g_type( Queue_7_io_deq_bits_payload_g_type )
  );
  Queue_7 Queue_8(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_8_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_enq_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_deq_ready( io_tiles_0_probe_ready ),
       .io_deq_valid( Queue_8_io_deq_valid ),
       .io_deq_bits_header_src( Queue_8_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_8_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_8_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_master_xact_id( Queue_8_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_p_type( Queue_8_io_deq_bits_payload_p_type )
  );
  Queue_3 Queue_9(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_9_io_enq_ready ),
       .io_enq_valid( T24 ),
       .io_enq_bits_header_src( T23 ),
       .io_enq_bits_header_dst( T22 ),
       .io_enq_bits_payload_addr( T21 ),
       .io_enq_bits_payload_client_xact_id( T20 ),
       .io_enq_bits_payload_data( T19 ),
       .io_enq_bits_payload_a_type( T18 ),
       .io_enq_bits_payload_write_mask( T17 ),
       .io_enq_bits_payload_subword_addr( T16 ),
       .io_enq_bits_payload_atomic_opcode( T15 ),
       .io_deq_ready( outmemsys_io_htif_acquire_ready ),
       .io_deq_valid( Queue_9_io_deq_valid ),
       .io_deq_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_9_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_9_io_deq_bits_payload_data ),
       .io_deq_bits_payload_a_type( Queue_9_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_write_mask( Queue_9_io_deq_bits_payload_write_mask ),
       .io_deq_bits_payload_subword_addr( Queue_9_io_deq_bits_payload_subword_addr ),
       .io_deq_bits_payload_atomic_opcode( Queue_9_io_deq_bits_payload_atomic_opcode )
  );
  Queue_4 Queue_10(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_10_io_enq_ready ),
       .io_enq_valid( T14 ),
       .io_enq_bits_header_src( T13 ),
       .io_enq_bits_header_dst( T12 ),
       .io_enq_bits_payload_addr( T11 ),
       .io_enq_bits_payload_client_xact_id( T10 ),
       .io_enq_bits_payload_master_xact_id( T9 ),
       .io_enq_bits_payload_data( T8 ),
       .io_enq_bits_payload_r_type( T7 ),
       .io_deq_ready( outmemsys_io_htif_release_ready ),
       .io_deq_valid( Queue_10_io_deq_valid ),
       .io_deq_bits_header_src( Queue_10_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_10_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_10_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_10_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_10_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_data( Queue_10_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_10_io_deq_bits_payload_r_type )
  );
  Queue_5 Queue_11(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_11_io_enq_ready ),
       .io_enq_valid( T6 ),
       .io_enq_bits_header_src( T5 ),
       .io_enq_bits_header_dst( T4 ),
       .io_enq_bits_payload_master_xact_id( T3 ),
       .io_deq_ready( outmemsys_io_htif_finish_ready ),
       .io_deq_valid( Queue_11_io_deq_valid ),
       .io_deq_bits_header_src( Queue_11_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_11_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_11_io_deq_bits_payload_master_xact_id )
  );
  Queue_6 Queue_12(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_12_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_deq_ready( htif_io_mem_grant_ready ),
       .io_deq_valid( Queue_12_io_deq_valid ),
       .io_deq_bits_header_src( Queue_12_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_12_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_12_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_12_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_12_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_g_type( Queue_12_io_deq_bits_payload_g_type )
  );
  Queue_7 Queue_13(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_13_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_htif_probe_bits_payload_master_xact_id ),
       .io_enq_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_deq_ready( htif_io_mem_probe_ready ),
       .io_deq_valid( Queue_13_io_deq_valid ),
       .io_deq_bits_header_src( Queue_13_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_13_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_13_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_master_xact_id( Queue_13_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_p_type( Queue_13_io_deq_bits_payload_p_type )
  );
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [4:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[4:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data
);

  wire[63:0] T0;
  wire[69:0] T1;
  reg [69:0] ram [1:0];
  wire[69:0] T2;
  wire[69:0] T3;
  wire[69:0] T4;
  wire[68:0] T5;
  wire do_enq;
  reg  R6;
  wire T19;
  wire T7;
  wire T8;
  reg  R9;
  wire T20;
  wire T10;
  wire T11;
  wire do_deq;
  wire[4:0] T12;
  wire T13;
  wire T14;
  wire empty;
  wire T15;
  reg  maybe_full;
  wire T21;
  wire T16;
  wire T17;
  wire ptr_match;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
    R6 = {1{$random}};
    R9 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[6'h3f:1'h0];
  assign T1 = ram[R9];
  assign T3 = T4;
  assign T4 = {io_enq_bits_rw, T5};
  assign T5 = {io_enq_bits_addr, io_enq_bits_data};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T19 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R6;
  assign T8 = R6 + 1'h1;
  assign T20 = reset ? 1'h0 : T10;
  assign T10 = do_deq ? T11 : R9;
  assign T11 = R9 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_addr = T12;
  assign T12 = T1[7'h44:7'h40];
  assign io_deq_bits_rw = T13;
  assign T13 = T1[7'h45:7'h45];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = ptr_match & T15;
  assign T15 = maybe_full ^ 1'h1;
  assign T21 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign ptr_match = R6 == R9;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T8;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else if(do_deq) begin
      R9 <= T11;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits
);

  wire[63:0] T0;
  reg [63:0] ram [1:0];
  wire[63:0] T1;
  wire do_enq;
  reg  R2;
  wire T13;
  wire T3;
  wire T4;
  reg  R5;
  wire T14;
  wire T6;
  wire T7;
  wire do_deq;
  wire T8;
  wire empty;
  wire T9;
  reg  maybe_full;
  wire T15;
  wire T10;
  wire T11;
  wire ptr_match;
  wire T12;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
    R2 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[R5];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T13 = reset ? 1'h0 : T3;
  assign T3 = do_enq ? T4 : R2;
  assign T4 = R2 + 1'h1;
  assign T14 = reset ? 1'h0 : T6;
  assign T6 = do_deq ? T7 : R5;
  assign T7 = R5 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T8;
  assign T8 = empty ^ 1'h1;
  assign empty = ptr_match & T9;
  assign T9 = maybe_full ^ 1'h1;
  assign T15 = reset ? 1'h0 : T10;
  assign T10 = T11 ? do_enq : maybe_full;
  assign T11 = do_enq != do_deq;
  assign ptr_match = R2 == R5;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R2] <= io_enq_bits;
    if(reset) begin
      R2 <= 1'h0;
    end else if(do_enq) begin
      R2 <= T4;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_deq) begin
      R5 <= T7;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T11) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits
);

  wire T0;
  reg [0:0] ram [1:0];
  wire T1;
  wire do_enq;
  reg  R2;
  wire T13;
  wire T3;
  wire T4;
  reg  R5;
  wire T14;
  wire T6;
  wire T7;
  wire do_deq;
  wire T8;
  wire empty;
  wire T9;
  reg  maybe_full;
  wire T15;
  wire T10;
  wire T11;
  wire ptr_match;
  wire T12;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R2 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[R5];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T13 = reset ? 1'h0 : T3;
  assign T3 = do_enq ? T4 : R2;
  assign T4 = R2 + 1'h1;
  assign T14 = reset ? 1'h0 : T6;
  assign T6 = do_deq ? T7 : R5;
  assign T7 = R5 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T8;
  assign T8 = empty ^ 1'h1;
  assign empty = ptr_match & T9;
  assign T9 = maybe_full ^ 1'h1;
  assign T15 = reset ? 1'h0 : T10;
  assign T10 = T11 ? do_enq : maybe_full;
  assign T11 = do_enq != do_deq;
  assign ptr_match = R2 == R5;
  assign io_enq_ready = T12;
  assign T12 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R2] <= io_enq_bits;
    if(reset) begin
      R2 <= 1'h0;
    end else if(do_enq) begin
      R2 <= T4;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_deq) begin
      R5 <= T7;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T11) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Top(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    input  io_mem_backup_en,
    output io_in_mem_ready,
    input  io_in_mem_valid,
    input  io_out_mem_ready,
    output io_out_mem_valid
);

  wire resetSigs_0;
  reg  R0;
  reg  R1;
  wire Queue_0_io_enq_ready;
  wire Queue_0_io_deq_valid;
  wire Queue_0_io_deq_bits_rw;
  wire[4:0] Queue_0_io_deq_bits_addr;
  wire[63:0] Queue_0_io_deq_bits_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire Queue_2_io_deq_bits;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire Queue_3_io_deq_bits;
  wire Tile_io_tilelink_acquire_valid;
  wire[1:0] Tile_io_tilelink_acquire_bits_header_src;
  wire[1:0] Tile_io_tilelink_acquire_bits_header_dst;
  wire[25:0] Tile_io_tilelink_acquire_bits_payload_addr;
  wire[1:0] Tile_io_tilelink_acquire_bits_payload_client_xact_id;
  wire[511:0] Tile_io_tilelink_acquire_bits_payload_data;
  wire[2:0] Tile_io_tilelink_acquire_bits_payload_a_type;
  wire[5:0] Tile_io_tilelink_acquire_bits_payload_write_mask;
  wire[2:0] Tile_io_tilelink_acquire_bits_payload_subword_addr;
  wire[3:0] Tile_io_tilelink_acquire_bits_payload_atomic_opcode;
  wire Tile_io_tilelink_grant_ready;
  wire Tile_io_tilelink_finish_valid;
  wire[1:0] Tile_io_tilelink_finish_bits_header_src;
  wire[1:0] Tile_io_tilelink_finish_bits_header_dst;
  wire[2:0] Tile_io_tilelink_finish_bits_payload_master_xact_id;
  wire Tile_io_tilelink_probe_ready;
  wire Tile_io_tilelink_release_valid;
  wire[1:0] Tile_io_tilelink_release_bits_header_src;
  wire[1:0] Tile_io_tilelink_release_bits_header_dst;
  wire[25:0] Tile_io_tilelink_release_bits_payload_addr;
  wire[1:0] Tile_io_tilelink_release_bits_payload_client_xact_id;
  wire[2:0] Tile_io_tilelink_release_bits_payload_master_xact_id;
  wire[511:0] Tile_io_tilelink_release_bits_payload_data;
  wire[2:0] Tile_io_tilelink_release_bits_payload_r_type;
  wire Tile_io_host_pcr_req_ready;
  wire Tile_io_host_pcr_rep_valid;
  wire[63:0] Tile_io_host_pcr_rep_bits;
  wire Tile_io_host_ipi_req_valid;
  wire Tile_io_host_ipi_req_bits;
  wire Tile_io_host_ipi_rep_ready;
  wire Tile_io_host_debug_stats_pcr;
  wire uncore_io_host_in_ready;
  wire uncore_io_host_out_valid;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_debug_stats_pcr;
  wire uncore_io_mem_req_cmd_valid;
  wire[25:0] uncore_io_mem_req_cmd_bits_addr;
  wire[4:0] uncore_io_mem_req_cmd_bits_tag;
  wire uncore_io_mem_req_cmd_bits_rw;
  wire uncore_io_mem_req_data_valid;
  wire[127:0] uncore_io_mem_req_data_bits_data;
  wire uncore_io_tiles_0_acquire_ready;
  wire uncore_io_tiles_0_grant_valid;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_src;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_dst;
  wire[511:0] uncore_io_tiles_0_grant_bits_payload_data;
  wire[1:0] uncore_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[2:0] uncore_io_tiles_0_grant_bits_payload_master_xact_id;
  wire[3:0] uncore_io_tiles_0_grant_bits_payload_g_type;
  wire uncore_io_tiles_0_finish_ready;
  wire uncore_io_tiles_0_probe_valid;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_src;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_dst;
  wire[25:0] uncore_io_tiles_0_probe_bits_payload_addr;
  wire[2:0] uncore_io_tiles_0_probe_bits_payload_master_xact_id;
  wire[1:0] uncore_io_tiles_0_probe_bits_payload_p_type;
  wire uncore_io_tiles_0_release_ready;
  wire uncore_io_htif_0_reset;
  wire uncore_io_htif_0_pcr_req_valid;
  wire uncore_io_htif_0_pcr_req_bits_rw;
  wire[4:0] uncore_io_htif_0_pcr_req_bits_addr;
  wire[63:0] uncore_io_htif_0_pcr_req_bits_data;
  wire uncore_io_htif_0_pcr_rep_ready;
  wire uncore_io_htif_0_ipi_req_ready;
  wire uncore_io_htif_0_ipi_rep_valid;
  wire uncore_io_htif_0_ipi_rep_bits;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
  end
`endif

  assign resetSigs_0 = uncore_io_htif_0_reset;
  assign io_mem_req_data_bits_data = uncore_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = uncore_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = uncore_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = uncore_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = uncore_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = uncore_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = uncore_io_host_debug_stats_pcr;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
  Tile Tile(.clk(clk), .reset(resetSigs_0),
       .io_tilelink_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tilelink_acquire_valid( Tile_io_tilelink_acquire_valid ),
       .io_tilelink_acquire_bits_header_src( Tile_io_tilelink_acquire_bits_header_src ),
       .io_tilelink_acquire_bits_header_dst( Tile_io_tilelink_acquire_bits_header_dst ),
       .io_tilelink_acquire_bits_payload_addr( Tile_io_tilelink_acquire_bits_payload_addr ),
       .io_tilelink_acquire_bits_payload_client_xact_id( Tile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tilelink_acquire_bits_payload_data( Tile_io_tilelink_acquire_bits_payload_data ),
       .io_tilelink_acquire_bits_payload_a_type( Tile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tilelink_acquire_bits_payload_write_mask( Tile_io_tilelink_acquire_bits_payload_write_mask ),
       .io_tilelink_acquire_bits_payload_subword_addr( Tile_io_tilelink_acquire_bits_payload_subword_addr ),
       .io_tilelink_acquire_bits_payload_atomic_opcode( Tile_io_tilelink_acquire_bits_payload_atomic_opcode ),
       .io_tilelink_grant_ready( Tile_io_tilelink_grant_ready ),
       .io_tilelink_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tilelink_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tilelink_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tilelink_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tilelink_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tilelink_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tilelink_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tilelink_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tilelink_finish_valid( Tile_io_tilelink_finish_valid ),
       .io_tilelink_finish_bits_header_src( Tile_io_tilelink_finish_bits_header_src ),
       .io_tilelink_finish_bits_header_dst( Tile_io_tilelink_finish_bits_header_dst ),
       .io_tilelink_finish_bits_payload_master_xact_id( Tile_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tilelink_probe_ready( Tile_io_tilelink_probe_ready ),
       .io_tilelink_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tilelink_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tilelink_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tilelink_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tilelink_probe_bits_payload_master_xact_id( uncore_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tilelink_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tilelink_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tilelink_release_valid( Tile_io_tilelink_release_valid ),
       .io_tilelink_release_bits_header_src( Tile_io_tilelink_release_bits_header_src ),
       .io_tilelink_release_bits_header_dst( Tile_io_tilelink_release_bits_header_dst ),
       .io_tilelink_release_bits_payload_addr( Tile_io_tilelink_release_bits_payload_addr ),
       .io_tilelink_release_bits_payload_client_xact_id( Tile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tilelink_release_bits_payload_master_xact_id( Tile_io_tilelink_release_bits_payload_master_xact_id ),
       .io_tilelink_release_bits_payload_data( Tile_io_tilelink_release_bits_payload_data ),
       .io_tilelink_release_bits_payload_r_type( Tile_io_tilelink_release_bits_payload_r_type ),
       .io_host_reset( R0 ),
       .io_host_id( 1'h0 ),
       .io_host_pcr_req_ready( Tile_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( Queue_0_io_deq_valid ),
       .io_host_pcr_req_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_host_pcr_req_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_host_pcr_req_bits_data( Queue_0_io_deq_bits_data ),
       .io_host_pcr_rep_ready( Queue_1_io_enq_ready ),
       .io_host_pcr_rep_valid( Tile_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( Tile_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( Queue_2_io_enq_ready ),
       .io_host_ipi_req_valid( Tile_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( Tile_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( Tile_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( Queue_3_io_deq_valid ),
       .io_host_ipi_rep_bits( Queue_3_io_deq_bits ),
       .io_host_debug_stats_pcr( Tile_io_host_debug_stats_pcr )
  );
  Uncore uncore(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       .io_host_debug_stats_pcr( uncore_io_host_debug_stats_pcr ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( uncore_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( uncore_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( uncore_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( uncore_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( uncore_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( uncore_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag ),
       .io_tiles_0_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( Tile_io_tilelink_acquire_valid ),
       .io_tiles_0_acquire_bits_header_src( Tile_io_tilelink_acquire_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( Tile_io_tilelink_acquire_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( Tile_io_tilelink_acquire_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( Tile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( Tile_io_tilelink_acquire_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_a_type( Tile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_write_mask( Tile_io_tilelink_acquire_bits_payload_write_mask ),
       .io_tiles_0_acquire_bits_payload_subword_addr( Tile_io_tilelink_acquire_bits_payload_subword_addr ),
       .io_tiles_0_acquire_bits_payload_atomic_opcode( Tile_io_tilelink_acquire_bits_payload_atomic_opcode ),
       .io_tiles_0_grant_ready( Tile_io_tilelink_grant_ready ),
       .io_tiles_0_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( Tile_io_tilelink_finish_valid ),
       .io_tiles_0_finish_bits_header_src( Tile_io_tilelink_finish_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( Tile_io_tilelink_finish_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( Tile_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( Tile_io_tilelink_probe_ready ),
       .io_tiles_0_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_master_xact_id( uncore_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tiles_0_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( Tile_io_tilelink_release_valid ),
       .io_tiles_0_release_bits_header_src( Tile_io_tilelink_release_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( Tile_io_tilelink_release_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( Tile_io_tilelink_release_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( Tile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_master_xact_id( Tile_io_tilelink_release_bits_payload_master_xact_id ),
       .io_tiles_0_release_bits_payload_data( Tile_io_tilelink_release_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( Tile_io_tilelink_release_bits_payload_r_type ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_pcr_req_ready( Queue_0_io_enq_ready ),
       .io_htif_0_pcr_req_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_htif_0_pcr_req_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_htif_0_pcr_req_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_htif_0_pcr_req_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_htif_0_pcr_rep_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_htif_0_pcr_rep_valid( Queue_1_io_deq_valid ),
       .io_htif_0_pcr_rep_bits( Queue_1_io_deq_bits ),
       .io_htif_0_ipi_req_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_htif_0_ipi_req_valid( Queue_2_io_deq_valid ),
       .io_htif_0_ipi_req_bits( Queue_2_io_deq_bits ),
       .io_htif_0_ipi_rep_ready( Queue_3_io_enq_ready ),
       .io_htif_0_ipi_rep_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_htif_0_ipi_rep_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_htif_0_debug_stats_pcr( Tile_io_host_debug_stats_pcr ),
       .io_incoherent_0( uncore_io_htif_0_reset )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
  `ifndef SYNTHESIS
    assign uncore.io_htif_0_ipi_rep_bits = {1{$random}};
  `endif
  Queue_0 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_deq_ready( Tile_io_host_pcr_req_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_0_io_deq_bits_data )
  );
  Queue_1 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( Tile_io_host_pcr_rep_valid ),
       .io_enq_bits( Tile_io_host_pcr_rep_bits ),
       .io_deq_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
  );
  Queue_2 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( Tile_io_host_ipi_req_valid ),
       .io_enq_bits( Tile_io_host_ipi_req_bits ),
       .io_deq_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits( Queue_2_io_deq_bits )
  );
  Queue_2 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_enq_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_deq_ready( Tile_io_host_ipi_rep_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits( Queue_3_io_deq_bits )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= uncore_io_htif_0_reset;
  end
endmodule

module DataArray_T1(
  input CLK,
  input RST,
  input init,
  input [7:0] W0A,
  input W0E,
  input [127:0] W0I,
  input [127:0] W0M,
  input [7:0] R1A,
  input R1E,
  output [127:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+64) begin
    for (j=1; j<64; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][63:0] <= W0I[63:0];
  if (W0E && W0M[64]) ram[W0A][127:64] <= W0I[127:64];
end
assign R1O = ram[reg_R1A];

endmodule


module MetadataArray_tag_arr(
  input CLK,
  input RST,
  input init,
  input [5:0] W0A,
  input W0E,
  input [21:0] W0I,
  input [21:0] W0M,
  input [5:0] R1A,
  input R1E,
  output [21:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<1; i=i+22) begin
    for (j=1; j<22; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [21:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [5:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][21:0] <= W0I[21:0];
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_tag_array(
  input CLK,
  input RST,
  input init,
  input [5:0] RW0A,
  input RW0E,
  input RW0W,
  input [19:0] RW0M,
  input [19:0] RW0I,
  output [19:0] RW0O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<1; i=i+20) begin
    for (j=1; j<20; j=j+1) begin
      if (RW0M[i] != RW0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [19:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [5:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W && RW0M[0]) ram[RW0A][19:0] <= RW0I[19:0];
end
assign RW0O = ram[reg_RW0A];

endmodule


module ICache_T103(
  input CLK,
  input RST,
  input init,
  input [7:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0I,
  output [127:0] RW0O
);

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W) ram[RW0A] <= RW0I;
end
assign RW0O = ram[reg_RW0A];

endmodule


module HellaFlowQueue_ram(
  input CLK,
  input RST,
  input init,
  input [4:0] W0A,
  input W0E,
  input [132:0] W0I,
  input [4:0] R1A,
  input R1E,
  output [132:0] R1O
);

reg [132:0] ram [31:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 32; initvar = initvar+1)
        ram[initvar] = {5 {$random}};
    end
  `endif
  reg [4:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


